/**************************************************************** 
  ** Title : on chip module
  ** Project :  full-search block matching algorithm on VLSI
***************************************************************** 
  ** File :  me_on_chip.v
  ** Author : fzp
  ** Organization: sjtu
  ** Created :  
  ** Last update : 
  ** Platform : 
  ** Simulators : 
  ** Synthesizers: 
  ** Targets : 
  ** Dependency :  
***************************************************************** 
  ** Description:  
***************************************************************** 
  ** Copyright (c) notice  
*****************************************************************/ 

//pin 
//32 data
//1 clk
//1 rst_n
//1 initial
//1 output


module me_on_chip
#(
    parameter WORD_WIDETH = 8
)
(
    input a,
    output reg b
);
endmodule