/**************************************************************** 
  ** Title : testbench
  ** Project :  full-search block matching algorithm on VLSI
***************************************************************** 
  ** File :  testbench.v
  ** Author : fzp
  ** Organization: sjtu
  ** Created :  
  ** Last update : 
  ** Platform : 
  ** Simulators : 
  ** Synthesizers: 
  ** Targets : 
  ** Dependency :  
***************************************************************** 
  ** Description:  
***************************************************************** 
  ** Copyright (c) notice  
*****************************************************************/ 
initial


module testbench
(
    input [21:0] count,
    output [33:0] data
);
	reg [33:0] mem[4194304:0];

endmodule