/**************************************************************** 
  ** Title : 19*19*8bit register
  ** Project :  full-search block matching algorithm on VLSI
***************************************************************** 
  ** File :  mem19198.v
  ** Author : fzp
  ** Organization: sjtu
  ** Created :  
  ** Last update : 
  ** Platform : 
  ** Simulators : 
  ** Synthesizers: 
  ** Targets : 
  ** Dependency :  
***************************************************************** 
  ** Description:  
***************************************************************** 
  ** Copyright (c) notice  
*****************************************************************/ 
module mem19198(
    input                       clk,
    input       [151:0]         buffer1,
    output reg  [7:0]           mem0000,
    output reg  [7:0]           mem0001,
    output reg  [7:0]           mem0002,
    output reg  [7:0]           mem0003,
    output reg  [7:0]           mem0004,
    output reg  [7:0]           mem0005,
    output reg  [7:0]           mem0006,
    output reg  [7:0]           mem0007,
    output reg  [7:0]           mem0008,
    output reg  [7:0]           mem0009,
    output reg  [7:0]           mem0010,
    output reg  [7:0]           mem0011,
    output reg  [7:0]           mem0012,
    output reg  [7:0]           mem0013,
    output reg  [7:0]           mem0014,
    output reg  [7:0]           mem0015,
    output reg  [7:0]           mem0016,
    output reg  [7:0]           mem0017,
    output reg  [7:0]           mem0018,
    output reg  [7:0]           mem0100,
    output reg  [7:0]           mem0101,
    output reg  [7:0]           mem0102,
    output reg  [7:0]           mem0103,
    output reg  [7:0]           mem0104,
    output reg  [7:0]           mem0105,
    output reg  [7:0]           mem0106,
    output reg  [7:0]           mem0107,
    output reg  [7:0]           mem0108,
    output reg  [7:0]           mem0109,
    output reg  [7:0]           mem0110,
    output reg  [7:0]           mem0111,
    output reg  [7:0]           mem0112,
    output reg  [7:0]           mem0113,
    output reg  [7:0]           mem0114,
    output reg  [7:0]           mem0115,
    output reg  [7:0]           mem0116,
    output reg  [7:0]           mem0117,
    output reg  [7:0]           mem0118,
    output reg  [7:0]           mem0200,
    output reg  [7:0]           mem0201,
    output reg  [7:0]           mem0202,
    output reg  [7:0]           mem0203,
    output reg  [7:0]           mem0204,
    output reg  [7:0]           mem0205,
    output reg  [7:0]           mem0206,
    output reg  [7:0]           mem0207,
    output reg  [7:0]           mem0208,
    output reg  [7:0]           mem0209,
    output reg  [7:0]           mem0210,
    output reg  [7:0]           mem0211,
    output reg  [7:0]           mem0212,
    output reg  [7:0]           mem0213,
    output reg  [7:0]           mem0214,
    output reg  [7:0]           mem0215,
    output reg  [7:0]           mem0216,
    output reg  [7:0]           mem0217,
    output reg  [7:0]           mem0218,
    output reg  [7:0]           mem0300,
    output reg  [7:0]           mem0301,
    output reg  [7:0]           mem0302,
    output reg  [7:0]           mem0303,
    output reg  [7:0]           mem0304,
    output reg  [7:0]           mem0305,
    output reg  [7:0]           mem0306,
    output reg  [7:0]           mem0307,
    output reg  [7:0]           mem0308,
    output reg  [7:0]           mem0309,
    output reg  [7:0]           mem0310,
    output reg  [7:0]           mem0311,
    output reg  [7:0]           mem0312,
    output reg  [7:0]           mem0313,
    output reg  [7:0]           mem0314,
    output reg  [7:0]           mem0315,
    output reg  [7:0]           mem0316,
    output reg  [7:0]           mem0317,
    output reg  [7:0]           mem0318,
    output reg  [7:0]           mem0400,
    output reg  [7:0]           mem0401,
    output reg  [7:0]           mem0402,
    output reg  [7:0]           mem0403,
    output reg  [7:0]           mem0404,
    output reg  [7:0]           mem0405,
    output reg  [7:0]           mem0406,
    output reg  [7:0]           mem0407,
    output reg  [7:0]           mem0408,
    output reg  [7:0]           mem0409,
    output reg  [7:0]           mem0410,
    output reg  [7:0]           mem0411,
    output reg  [7:0]           mem0412,
    output reg  [7:0]           mem0413,
    output reg  [7:0]           mem0414,
    output reg  [7:0]           mem0415,
    output reg  [7:0]           mem0416,
    output reg  [7:0]           mem0417,
    output reg  [7:0]           mem0418,
    output reg  [7:0]           mem0500,
    output reg  [7:0]           mem0501,
    output reg  [7:0]           mem0502,
    output reg  [7:0]           mem0503,
    output reg  [7:0]           mem0504,
    output reg  [7:0]           mem0505,
    output reg  [7:0]           mem0506,
    output reg  [7:0]           mem0507,
    output reg  [7:0]           mem0508,
    output reg  [7:0]           mem0509,
    output reg  [7:0]           mem0510,
    output reg  [7:0]           mem0511,
    output reg  [7:0]           mem0512,
    output reg  [7:0]           mem0513,
    output reg  [7:0]           mem0514,
    output reg  [7:0]           mem0515,
    output reg  [7:0]           mem0516,
    output reg  [7:0]           mem0517,
    output reg  [7:0]           mem0518,
    output reg  [7:0]           mem0600,
    output reg  [7:0]           mem0601,
    output reg  [7:0]           mem0602,
    output reg  [7:0]           mem0603,
    output reg  [7:0]           mem0604,
    output reg  [7:0]           mem0605,
    output reg  [7:0]           mem0606,
    output reg  [7:0]           mem0607,
    output reg  [7:0]           mem0608,
    output reg  [7:0]           mem0609,
    output reg  [7:0]           mem0610,
    output reg  [7:0]           mem0611,
    output reg  [7:0]           mem0612,
    output reg  [7:0]           mem0613,
    output reg  [7:0]           mem0614,
    output reg  [7:0]           mem0615,
    output reg  [7:0]           mem0616,
    output reg  [7:0]           mem0617,
    output reg  [7:0]           mem0618,
    output reg  [7:0]           mem0700,
    output reg  [7:0]           mem0701,
    output reg  [7:0]           mem0702,
    output reg  [7:0]           mem0703,
    output reg  [7:0]           mem0704,
    output reg  [7:0]           mem0705,
    output reg  [7:0]           mem0706,
    output reg  [7:0]           mem0707,
    output reg  [7:0]           mem0708,
    output reg  [7:0]           mem0709,
    output reg  [7:0]           mem0710,
    output reg  [7:0]           mem0711,
    output reg  [7:0]           mem0712,
    output reg  [7:0]           mem0713,
    output reg  [7:0]           mem0714,
    output reg  [7:0]           mem0715,
    output reg  [7:0]           mem0716,
    output reg  [7:0]           mem0717,
    output reg  [7:0]           mem0718,
    output reg  [7:0]           mem0800,
    output reg  [7:0]           mem0801,
    output reg  [7:0]           mem0802,
    output reg  [7:0]           mem0803,
    output reg  [7:0]           mem0804,
    output reg  [7:0]           mem0805,
    output reg  [7:0]           mem0806,
    output reg  [7:0]           mem0807,
    output reg  [7:0]           mem0808,
    output reg  [7:0]           mem0809,
    output reg  [7:0]           mem0810,
    output reg  [7:0]           mem0811,
    output reg  [7:0]           mem0812,
    output reg  [7:0]           mem0813,
    output reg  [7:0]           mem0814,
    output reg  [7:0]           mem0815,
    output reg  [7:0]           mem0816,
    output reg  [7:0]           mem0817,
    output reg  [7:0]           mem0818,
    output reg  [7:0]           mem0900,
    output reg  [7:0]           mem0901,
    output reg  [7:0]           mem0902,
    output reg  [7:0]           mem0903,
    output reg  [7:0]           mem0904,
    output reg  [7:0]           mem0905,
    output reg  [7:0]           mem0906,
    output reg  [7:0]           mem0907,
    output reg  [7:0]           mem0908,
    output reg  [7:0]           mem0909,
    output reg  [7:0]           mem0910,
    output reg  [7:0]           mem0911,
    output reg  [7:0]           mem0912,
    output reg  [7:0]           mem0913,
    output reg  [7:0]           mem0914,
    output reg  [7:0]           mem0915,
    output reg  [7:0]           mem0916,
    output reg  [7:0]           mem0917,
    output reg  [7:0]           mem0918,
    output reg  [7:0]           mem1000,
    output reg  [7:0]           mem1001,
    output reg  [7:0]           mem1002,
    output reg  [7:0]           mem1003,
    output reg  [7:0]           mem1004,
    output reg  [7:0]           mem1005,
    output reg  [7:0]           mem1006,
    output reg  [7:0]           mem1007,
    output reg  [7:0]           mem1008,
    output reg  [7:0]           mem1009,
    output reg  [7:0]           mem1010,
    output reg  [7:0]           mem1011,
    output reg  [7:0]           mem1012,
    output reg  [7:0]           mem1013,
    output reg  [7:0]           mem1014,
    output reg  [7:0]           mem1015,
    output reg  [7:0]           mem1016,
    output reg  [7:0]           mem1017,
    output reg  [7:0]           mem1018,
    output reg  [7:0]           mem1100,
    output reg  [7:0]           mem1101,
    output reg  [7:0]           mem1102,
    output reg  [7:0]           mem1103,
    output reg  [7:0]           mem1104,
    output reg  [7:0]           mem1105,
    output reg  [7:0]           mem1106,
    output reg  [7:0]           mem1107,
    output reg  [7:0]           mem1108,
    output reg  [7:0]           mem1109,
    output reg  [7:0]           mem1110,
    output reg  [7:0]           mem1111,
    output reg  [7:0]           mem1112,
    output reg  [7:0]           mem1113,
    output reg  [7:0]           mem1114,
    output reg  [7:0]           mem1115,
    output reg  [7:0]           mem1116,
    output reg  [7:0]           mem1117,
    output reg  [7:0]           mem1118,
    output reg  [7:0]           mem1200,
    output reg  [7:0]           mem1201,
    output reg  [7:0]           mem1202,
    output reg  [7:0]           mem1203,
    output reg  [7:0]           mem1204,
    output reg  [7:0]           mem1205,
    output reg  [7:0]           mem1206,
    output reg  [7:0]           mem1207,
    output reg  [7:0]           mem1208,
    output reg  [7:0]           mem1209,
    output reg  [7:0]           mem1210,
    output reg  [7:0]           mem1211,
    output reg  [7:0]           mem1212,
    output reg  [7:0]           mem1213,
    output reg  [7:0]           mem1214,
    output reg  [7:0]           mem1215,
    output reg  [7:0]           mem1216,
    output reg  [7:0]           mem1217,
    output reg  [7:0]           mem1218,
    output reg  [7:0]           mem1300,
    output reg  [7:0]           mem1301,
    output reg  [7:0]           mem1302,
    output reg  [7:0]           mem1303,
    output reg  [7:0]           mem1304,
    output reg  [7:0]           mem1305,
    output reg  [7:0]           mem1306,
    output reg  [7:0]           mem1307,
    output reg  [7:0]           mem1308,
    output reg  [7:0]           mem1309,
    output reg  [7:0]           mem1310,
    output reg  [7:0]           mem1311,
    output reg  [7:0]           mem1312,
    output reg  [7:0]           mem1313,
    output reg  [7:0]           mem1314,
    output reg  [7:0]           mem1315,
    output reg  [7:0]           mem1316,
    output reg  [7:0]           mem1317,
    output reg  [7:0]           mem1318,
    output reg  [7:0]           mem1400,
    output reg  [7:0]           mem1401,
    output reg  [7:0]           mem1402,
    output reg  [7:0]           mem1403,
    output reg  [7:0]           mem1404,
    output reg  [7:0]           mem1405,
    output reg  [7:0]           mem1406,
    output reg  [7:0]           mem1407,
    output reg  [7:0]           mem1408,
    output reg  [7:0]           mem1409,
    output reg  [7:0]           mem1410,
    output reg  [7:0]           mem1411,
    output reg  [7:0]           mem1412,
    output reg  [7:0]           mem1413,
    output reg  [7:0]           mem1414,
    output reg  [7:0]           mem1415,
    output reg  [7:0]           mem1416,
    output reg  [7:0]           mem1417,
    output reg  [7:0]           mem1418,
    output reg  [7:0]           mem1500,
    output reg  [7:0]           mem1501,
    output reg  [7:0]           mem1502,
    output reg  [7:0]           mem1503,
    output reg  [7:0]           mem1504,
    output reg  [7:0]           mem1505,
    output reg  [7:0]           mem1506,
    output reg  [7:0]           mem1507,
    output reg  [7:0]           mem1508,
    output reg  [7:0]           mem1509,
    output reg  [7:0]           mem1510,
    output reg  [7:0]           mem1511,
    output reg  [7:0]           mem1512,
    output reg  [7:0]           mem1513,
    output reg  [7:0]           mem1514,
    output reg  [7:0]           mem1515,
    output reg  [7:0]           mem1516,
    output reg  [7:0]           mem1517,
    output reg  [7:0]           mem1518,
    output reg  [7:0]           mem1600,
    output reg  [7:0]           mem1601,
    output reg  [7:0]           mem1602,
    output reg  [7:0]           mem1603,
    output reg  [7:0]           mem1604,
    output reg  [7:0]           mem1605,
    output reg  [7:0]           mem1606,
    output reg  [7:0]           mem1607,
    output reg  [7:0]           mem1608,
    output reg  [7:0]           mem1609,
    output reg  [7:0]           mem1610,
    output reg  [7:0]           mem1611,
    output reg  [7:0]           mem1612,
    output reg  [7:0]           mem1613,
    output reg  [7:0]           mem1614,
    output reg  [7:0]           mem1615,
    output reg  [7:0]           mem1616,
    output reg  [7:0]           mem1617,
    output reg  [7:0]           mem1618,
    output reg  [7:0]           mem1700,
    output reg  [7:0]           mem1701,
    output reg  [7:0]           mem1702,
    output reg  [7:0]           mem1703,
    output reg  [7:0]           mem1704,
    output reg  [7:0]           mem1705,
    output reg  [7:0]           mem1706,
    output reg  [7:0]           mem1707,
    output reg  [7:0]           mem1708,
    output reg  [7:0]           mem1709,
    output reg  [7:0]           mem1710,
    output reg  [7:0]           mem1711,
    output reg  [7:0]           mem1712,
    output reg  [7:0]           mem1713,
    output reg  [7:0]           mem1714,
    output reg  [7:0]           mem1715,
    output reg  [7:0]           mem1716,
    output reg  [7:0]           mem1717,
    output reg  [7:0]           mem1718,
    output reg  [7:0]           mem1800,
    output reg  [7:0]           mem1801,
    output reg  [7:0]           mem1802,
    output reg  [7:0]           mem1803,
    output reg  [7:0]           mem1804,
    output reg  [7:0]           mem1805,
    output reg  [7:0]           mem1806,
    output reg  [7:0]           mem1807,
    output reg  [7:0]           mem1808,
    output reg  [7:0]           mem1809,
    output reg  [7:0]           mem1810,
    output reg  [7:0]           mem1811,
    output reg  [7:0]           mem1812,
    output reg  [7:0]           mem1813,
    output reg  [7:0]           mem1814,
    output reg  [7:0]           mem1815,
    output reg  [7:0]           mem1816,
    output reg  [7:0]           mem1817,
    output reg  [7:0]           mem1818
)

always @ (clk)
begin
  
end

endmodule