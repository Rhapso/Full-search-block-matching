/**************************************************************** 
  ** Title : 19*19*8bit register
  ** Project :  full-search block matching algorithm on VLSI
***************************************************************** 
  ** File :  mem19198.v
  ** Author : fzp
  ** Organization: sjtu
  ** Created :  
  ** Last update : 
  ** Platform : 
  ** Simulators : 
  ** Synthesizers: 
  ** Targets : 
  ** Dependency :  
***************************************************************** 
  ** Description:  
***************************************************************** 
  ** Copyright (c) notice  
*****************************************************************/ 


module mem19198
#(
    parameter   WORD_WIDETH         8,
    parameter   INPUT_DATA_PIN      32
)
(
    input                                   clk,
    input       [INPUT_DATA_PIN-1:0]        input_raw,
    input       [3:0]                       ctr_word,
    input                                   en_input,
    output reg  [WORD_WIDETH-1:0]           pe00_in00,
    output reg  [WORD_WIDETH-1:0]           pe00_in01,
    output reg  [WORD_WIDETH-1:0]           pe00_in02,
    output reg  [WORD_WIDETH-1:0]           pe00_in03,
    output reg  [WORD_WIDETH-1:0]           pe00_in04,
    output reg  [WORD_WIDETH-1:0]           pe00_in05,
    output reg  [WORD_WIDETH-1:0]           pe00_in06,
    output reg  [WORD_WIDETH-1:0]           pe00_in07,
    output reg  [WORD_WIDETH-1:0]           pe00_in08,
    output reg  [WORD_WIDETH-1:0]           pe00_in09,
    output reg  [WORD_WIDETH-1:0]           pe00_in10,
    output reg  [WORD_WIDETH-1:0]           pe00_in11,
    output reg  [WORD_WIDETH-1:0]           pe00_in12,
    output reg  [WORD_WIDETH-1:0]           pe00_in13,
    output reg  [WORD_WIDETH-1:0]           pe00_in14,
    output reg  [WORD_WIDETH-1:0]           pe00_in15,
    output reg  [WORD_WIDETH-1:0]           pe01_in00,
    output reg  [WORD_WIDETH-1:0]           pe01_in01,
    output reg  [WORD_WIDETH-1:0]           pe01_in02,
    output reg  [WORD_WIDETH-1:0]           pe01_in03,
    output reg  [WORD_WIDETH-1:0]           pe01_in04,
    output reg  [WORD_WIDETH-1:0]           pe01_in05,
    output reg  [WORD_WIDETH-1:0]           pe01_in06,
    output reg  [WORD_WIDETH-1:0]           pe01_in07,
    output reg  [WORD_WIDETH-1:0]           pe01_in08,
    output reg  [WORD_WIDETH-1:0]           pe01_in09,
    output reg  [WORD_WIDETH-1:0]           pe01_in10,
    output reg  [WORD_WIDETH-1:0]           pe01_in11,
    output reg  [WORD_WIDETH-1:0]           pe01_in12,
    output reg  [WORD_WIDETH-1:0]           pe01_in13,
    output reg  [WORD_WIDETH-1:0]           pe01_in14,
    output reg  [WORD_WIDETH-1:0]           pe01_in15,
    output reg  [WORD_WIDETH-1:0]           pe02_in00,
    output reg  [WORD_WIDETH-1:0]           pe02_in01,
    output reg  [WORD_WIDETH-1:0]           pe02_in02,
    output reg  [WORD_WIDETH-1:0]           pe02_in03,
    output reg  [WORD_WIDETH-1:0]           pe02_in04,
    output reg  [WORD_WIDETH-1:0]           pe02_in05,
    output reg  [WORD_WIDETH-1:0]           pe02_in06,
    output reg  [WORD_WIDETH-1:0]           pe02_in07,
    output reg  [WORD_WIDETH-1:0]           pe02_in08,
    output reg  [WORD_WIDETH-1:0]           pe02_in09,
    output reg  [WORD_WIDETH-1:0]           pe02_in10,
    output reg  [WORD_WIDETH-1:0]           pe02_in11,
    output reg  [WORD_WIDETH-1:0]           pe02_in12,
    output reg  [WORD_WIDETH-1:0]           pe02_in13,
    output reg  [WORD_WIDETH-1:0]           pe02_in14,
    output reg  [WORD_WIDETH-1:0]           pe02_in15,
    output reg  [WORD_WIDETH-1:0]           pe03_in00,
    output reg  [WORD_WIDETH-1:0]           pe03_in01,
    output reg  [WORD_WIDETH-1:0]           pe03_in02,
    output reg  [WORD_WIDETH-1:0]           pe03_in03,
    output reg  [WORD_WIDETH-1:0]           pe03_in04,
    output reg  [WORD_WIDETH-1:0]           pe03_in05,
    output reg  [WORD_WIDETH-1:0]           pe03_in06,
    output reg  [WORD_WIDETH-1:0]           pe03_in07,
    output reg  [WORD_WIDETH-1:0]           pe03_in08,
    output reg  [WORD_WIDETH-1:0]           pe03_in09,
    output reg  [WORD_WIDETH-1:0]           pe03_in10,
    output reg  [WORD_WIDETH-1:0]           pe03_in11,
    output reg  [WORD_WIDETH-1:0]           pe03_in12,
    output reg  [WORD_WIDETH-1:0]           pe03_in13,
    output reg  [WORD_WIDETH-1:0]           pe03_in14,
    output reg  [WORD_WIDETH-1:0]           pe03_in15,
    output reg  [WORD_WIDETH-1:0]           pe04_in00,
    output reg  [WORD_WIDETH-1:0]           pe04_in01,
    output reg  [WORD_WIDETH-1:0]           pe04_in02,
    output reg  [WORD_WIDETH-1:0]           pe04_in03,
    output reg  [WORD_WIDETH-1:0]           pe04_in04,
    output reg  [WORD_WIDETH-1:0]           pe04_in05,
    output reg  [WORD_WIDETH-1:0]           pe04_in06,
    output reg  [WORD_WIDETH-1:0]           pe04_in07,
    output reg  [WORD_WIDETH-1:0]           pe04_in08,
    output reg  [WORD_WIDETH-1:0]           pe04_in09,
    output reg  [WORD_WIDETH-1:0]           pe04_in10,
    output reg  [WORD_WIDETH-1:0]           pe04_in11,
    output reg  [WORD_WIDETH-1:0]           pe04_in12,
    output reg  [WORD_WIDETH-1:0]           pe04_in13,
    output reg  [WORD_WIDETH-1:0]           pe04_in14,
    output reg  [WORD_WIDETH-1:0]           pe04_in15,
    output reg  [WORD_WIDETH-1:0]           pe05_in00,
    output reg  [WORD_WIDETH-1:0]           pe05_in01,
    output reg  [WORD_WIDETH-1:0]           pe05_in02,
    output reg  [WORD_WIDETH-1:0]           pe05_in03,
    output reg  [WORD_WIDETH-1:0]           pe05_in04,
    output reg  [WORD_WIDETH-1:0]           pe05_in05,
    output reg  [WORD_WIDETH-1:0]           pe05_in06,
    output reg  [WORD_WIDETH-1:0]           pe05_in07,
    output reg  [WORD_WIDETH-1:0]           pe05_in08,
    output reg  [WORD_WIDETH-1:0]           pe05_in09,
    output reg  [WORD_WIDETH-1:0]           pe05_in10,
    output reg  [WORD_WIDETH-1:0]           pe05_in11,
    output reg  [WORD_WIDETH-1:0]           pe05_in12,
    output reg  [WORD_WIDETH-1:0]           pe05_in13,
    output reg  [WORD_WIDETH-1:0]           pe05_in14,
    output reg  [WORD_WIDETH-1:0]           pe05_in15,
    output reg  [WORD_WIDETH-1:0]           pe06_in00,
    output reg  [WORD_WIDETH-1:0]           pe06_in01,
    output reg  [WORD_WIDETH-1:0]           pe06_in02,
    output reg  [WORD_WIDETH-1:0]           pe06_in03,
    output reg  [WORD_WIDETH-1:0]           pe06_in04,
    output reg  [WORD_WIDETH-1:0]           pe06_in05,
    output reg  [WORD_WIDETH-1:0]           pe06_in06,
    output reg  [WORD_WIDETH-1:0]           pe06_in07,
    output reg  [WORD_WIDETH-1:0]           pe06_in08,
    output reg  [WORD_WIDETH-1:0]           pe06_in09,
    output reg  [WORD_WIDETH-1:0]           pe06_in10,
    output reg  [WORD_WIDETH-1:0]           pe06_in11,
    output reg  [WORD_WIDETH-1:0]           pe06_in12,
    output reg  [WORD_WIDETH-1:0]           pe06_in13,
    output reg  [WORD_WIDETH-1:0]           pe06_in14,
    output reg  [WORD_WIDETH-1:0]           pe06_in15,
    output reg  [WORD_WIDETH-1:0]           pe07_in00,
    output reg  [WORD_WIDETH-1:0]           pe07_in01,
    output reg  [WORD_WIDETH-1:0]           pe07_in02,
    output reg  [WORD_WIDETH-1:0]           pe07_in03,
    output reg  [WORD_WIDETH-1:0]           pe07_in04,
    output reg  [WORD_WIDETH-1:0]           pe07_in05,
    output reg  [WORD_WIDETH-1:0]           pe07_in06,
    output reg  [WORD_WIDETH-1:0]           pe07_in07,
    output reg  [WORD_WIDETH-1:0]           pe07_in08,
    output reg  [WORD_WIDETH-1:0]           pe07_in09,
    output reg  [WORD_WIDETH-1:0]           pe07_in10,
    output reg  [WORD_WIDETH-1:0]           pe07_in11,
    output reg  [WORD_WIDETH-1:0]           pe07_in12,
    output reg  [WORD_WIDETH-1:0]           pe07_in13,
    output reg  [WORD_WIDETH-1:0]           pe07_in14,
    output reg  [WORD_WIDETH-1:0]           pe07_in15,
    output reg  [WORD_WIDETH-1:0]           pe08_in00,
    output reg  [WORD_WIDETH-1:0]           pe08_in01,
    output reg  [WORD_WIDETH-1:0]           pe08_in02,
    output reg  [WORD_WIDETH-1:0]           pe08_in03,
    output reg  [WORD_WIDETH-1:0]           pe08_in04,
    output reg  [WORD_WIDETH-1:0]           pe08_in05,
    output reg  [WORD_WIDETH-1:0]           pe08_in06,
    output reg  [WORD_WIDETH-1:0]           pe08_in07,
    output reg  [WORD_WIDETH-1:0]           pe08_in08,
    output reg  [WORD_WIDETH-1:0]           pe08_in09,
    output reg  [WORD_WIDETH-1:0]           pe08_in10,
    output reg  [WORD_WIDETH-1:0]           pe08_in11,
    output reg  [WORD_WIDETH-1:0]           pe08_in12,
    output reg  [WORD_WIDETH-1:0]           pe08_in13,
    output reg  [WORD_WIDETH-1:0]           pe08_in14,
    output reg  [WORD_WIDETH-1:0]           pe08_in15,
    output reg  [WORD_WIDETH-1:0]           pe09_in00,
    output reg  [WORD_WIDETH-1:0]           pe09_in01,
    output reg  [WORD_WIDETH-1:0]           pe09_in02,
    output reg  [WORD_WIDETH-1:0]           pe09_in03,
    output reg  [WORD_WIDETH-1:0]           pe09_in04,
    output reg  [WORD_WIDETH-1:0]           pe09_in05,
    output reg  [WORD_WIDETH-1:0]           pe09_in06,
    output reg  [WORD_WIDETH-1:0]           pe09_in07,
    output reg  [WORD_WIDETH-1:0]           pe09_in08,
    output reg  [WORD_WIDETH-1:0]           pe09_in09,
    output reg  [WORD_WIDETH-1:0]           pe09_in10,
    output reg  [WORD_WIDETH-1:0]           pe09_in11,
    output reg  [WORD_WIDETH-1:0]           pe09_in12,
    output reg  [WORD_WIDETH-1:0]           pe09_in13,
    output reg  [WORD_WIDETH-1:0]           pe09_in14,
    output reg  [WORD_WIDETH-1:0]           pe09_in15,
    output reg  [WORD_WIDETH-1:0]           pe10_in00,
    output reg  [WORD_WIDETH-1:0]           pe10_in01,
    output reg  [WORD_WIDETH-1:0]           pe10_in02,
    output reg  [WORD_WIDETH-1:0]           pe10_in03,
    output reg  [WORD_WIDETH-1:0]           pe10_in04,
    output reg  [WORD_WIDETH-1:0]           pe10_in05,
    output reg  [WORD_WIDETH-1:0]           pe10_in06,
    output reg  [WORD_WIDETH-1:0]           pe10_in07,
    output reg  [WORD_WIDETH-1:0]           pe10_in08,
    output reg  [WORD_WIDETH-1:0]           pe10_in09,
    output reg  [WORD_WIDETH-1:0]           pe10_in10,
    output reg  [WORD_WIDETH-1:0]           pe10_in11,
    output reg  [WORD_WIDETH-1:0]           pe10_in12,
    output reg  [WORD_WIDETH-1:0]           pe10_in13,
    output reg  [WORD_WIDETH-1:0]           pe10_in14,
    output reg  [WORD_WIDETH-1:0]           pe10_in15,
    output reg  [WORD_WIDETH-1:0]           pe11_in00,
    output reg  [WORD_WIDETH-1:0]           pe11_in01,
    output reg  [WORD_WIDETH-1:0]           pe11_in02,
    output reg  [WORD_WIDETH-1:0]           pe11_in03,
    output reg  [WORD_WIDETH-1:0]           pe11_in04,
    output reg  [WORD_WIDETH-1:0]           pe11_in05,
    output reg  [WORD_WIDETH-1:0]           pe11_in06,
    output reg  [WORD_WIDETH-1:0]           pe11_in07,
    output reg  [WORD_WIDETH-1:0]           pe11_in08,
    output reg  [WORD_WIDETH-1:0]           pe11_in09,
    output reg  [WORD_WIDETH-1:0]           pe11_in10,
    output reg  [WORD_WIDETH-1:0]           pe11_in11,
    output reg  [WORD_WIDETH-1:0]           pe11_in12,
    output reg  [WORD_WIDETH-1:0]           pe11_in13,
    output reg  [WORD_WIDETH-1:0]           pe11_in14,
    output reg  [WORD_WIDETH-1:0]           pe11_in15,
    output reg  [WORD_WIDETH-1:0]           pe12_in00,
    output reg  [WORD_WIDETH-1:0]           pe12_in01,
    output reg  [WORD_WIDETH-1:0]           pe12_in02,
    output reg  [WORD_WIDETH-1:0]           pe12_in03,
    output reg  [WORD_WIDETH-1:0]           pe12_in04,
    output reg  [WORD_WIDETH-1:0]           pe12_in05,
    output reg  [WORD_WIDETH-1:0]           pe12_in06,
    output reg  [WORD_WIDETH-1:0]           pe12_in07,
    output reg  [WORD_WIDETH-1:0]           pe12_in08,
    output reg  [WORD_WIDETH-1:0]           pe12_in09,
    output reg  [WORD_WIDETH-1:0]           pe12_in10,
    output reg  [WORD_WIDETH-1:0]           pe12_in11,
    output reg  [WORD_WIDETH-1:0]           pe12_in12,
    output reg  [WORD_WIDETH-1:0]           pe12_in13,
    output reg  [WORD_WIDETH-1:0]           pe12_in14,
    output reg  [WORD_WIDETH-1:0]           pe12_in15,
    output reg  [WORD_WIDETH-1:0]           pe13_in00,
    output reg  [WORD_WIDETH-1:0]           pe13_in01,
    output reg  [WORD_WIDETH-1:0]           pe13_in02,
    output reg  [WORD_WIDETH-1:0]           pe13_in03,
    output reg  [WORD_WIDETH-1:0]           pe13_in04,
    output reg  [WORD_WIDETH-1:0]           pe13_in05,
    output reg  [WORD_WIDETH-1:0]           pe13_in06,
    output reg  [WORD_WIDETH-1:0]           pe13_in07,
    output reg  [WORD_WIDETH-1:0]           pe13_in08,
    output reg  [WORD_WIDETH-1:0]           pe13_in09,
    output reg  [WORD_WIDETH-1:0]           pe13_in10,
    output reg  [WORD_WIDETH-1:0]           pe13_in11,
    output reg  [WORD_WIDETH-1:0]           pe13_in12,
    output reg  [WORD_WIDETH-1:0]           pe13_in13,
    output reg  [WORD_WIDETH-1:0]           pe13_in14,
    output reg  [WORD_WIDETH-1:0]           pe13_in15,
    output reg  [WORD_WIDETH-1:0]           pe14_in00,
    output reg  [WORD_WIDETH-1:0]           pe14_in01,
    output reg  [WORD_WIDETH-1:0]           pe14_in02,
    output reg  [WORD_WIDETH-1:0]           pe14_in03,
    output reg  [WORD_WIDETH-1:0]           pe14_in04,
    output reg  [WORD_WIDETH-1:0]           pe14_in05,
    output reg  [WORD_WIDETH-1:0]           pe14_in06,
    output reg  [WORD_WIDETH-1:0]           pe14_in07,
    output reg  [WORD_WIDETH-1:0]           pe14_in08,
    output reg  [WORD_WIDETH-1:0]           pe14_in09,
    output reg  [WORD_WIDETH-1:0]           pe14_in10,
    output reg  [WORD_WIDETH-1:0]           pe14_in11,
    output reg  [WORD_WIDETH-1:0]           pe14_in12,
    output reg  [WORD_WIDETH-1:0]           pe14_in13,
    output reg  [WORD_WIDETH-1:0]           pe14_in14,
    output reg  [WORD_WIDETH-1:0]           pe14_in15,
    output reg  [WORD_WIDETH-1:0]           pe15_in00,
    output reg  [WORD_WIDETH-1:0]           pe15_in01,
    output reg  [WORD_WIDETH-1:0]           pe15_in02,
    output reg  [WORD_WIDETH-1:0]           pe15_in03,
    output reg  [WORD_WIDETH-1:0]           pe15_in04,
    output reg  [WORD_WIDETH-1:0]           pe15_in05,
    output reg  [WORD_WIDETH-1:0]           pe15_in06,
    output reg  [WORD_WIDETH-1:0]           pe15_in07,
    output reg  [WORD_WIDETH-1:0]           pe15_in08,
    output reg  [WORD_WIDETH-1:0]           pe15_in09,
    output reg  [WORD_WIDETH-1:0]           pe15_in10,
    output reg  [WORD_WIDETH-1:0]           pe15_in11,
    output reg  [WORD_WIDETH-1:0]           pe15_in12,
    output reg  [WORD_WIDETH-1:0]           pe15_in13,
    output reg  [WORD_WIDETH-1:0]           pe15_in14,
    output reg  [WORD_WIDETH-1:0]           pe15_in15
);
reg [WORD_WIDETH-1:0]           mem0000;
reg [WORD_WIDETH-1:0]           mem0001;
reg [WORD_WIDETH-1:0]           mem0002;
reg [WORD_WIDETH-1:0]           mem0003;
reg [WORD_WIDETH-1:0]           mem0004;
reg [WORD_WIDETH-1:0]           mem0005;
reg [WORD_WIDETH-1:0]           mem0006;
reg [WORD_WIDETH-1:0]           mem0007;
reg [WORD_WIDETH-1:0]           mem0008;
reg [WORD_WIDETH-1:0]           mem0009;
reg [WORD_WIDETH-1:0]           mem0010;
reg [WORD_WIDETH-1:0]           mem0011;
reg [WORD_WIDETH-1:0]           mem0012;
reg [WORD_WIDETH-1:0]           mem0013;
reg [WORD_WIDETH-1:0]           mem0014;
reg [WORD_WIDETH-1:0]           mem0015;
reg [WORD_WIDETH-1:0]           mem0016;
reg [WORD_WIDETH-1:0]           mem0017;
reg [WORD_WIDETH-1:0]           mem0018;
reg [WORD_WIDETH-1:0]           mem0100;
reg [WORD_WIDETH-1:0]           mem0101;
reg [WORD_WIDETH-1:0]           mem0102;
reg [WORD_WIDETH-1:0]           mem0103;
reg [WORD_WIDETH-1:0]           mem0104;
reg [WORD_WIDETH-1:0]           mem0105;
reg [WORD_WIDETH-1:0]           mem0106;
reg [WORD_WIDETH-1:0]           mem0107;
reg [WORD_WIDETH-1:0]           mem0108;
reg [WORD_WIDETH-1:0]           mem0109;
reg [WORD_WIDETH-1:0]           mem0110;
reg [WORD_WIDETH-1:0]           mem0111;
reg [WORD_WIDETH-1:0]           mem0112;
reg [WORD_WIDETH-1:0]           mem0113;
reg [WORD_WIDETH-1:0]           mem0114;
reg [WORD_WIDETH-1:0]           mem0115;
reg [WORD_WIDETH-1:0]           mem0116;
reg [WORD_WIDETH-1:0]           mem0117;
reg [WORD_WIDETH-1:0]           mem0118;
reg [WORD_WIDETH-1:0]           mem0200;
reg [WORD_WIDETH-1:0]           mem0201;
reg [WORD_WIDETH-1:0]           mem0202;
reg [WORD_WIDETH-1:0]           mem0203;
reg [WORD_WIDETH-1:0]           mem0204;
reg [WORD_WIDETH-1:0]           mem0205;
reg [WORD_WIDETH-1:0]           mem0206;
reg [WORD_WIDETH-1:0]           mem0207;
reg [WORD_WIDETH-1:0]           mem0208;
reg [WORD_WIDETH-1:0]           mem0209;
reg [WORD_WIDETH-1:0]           mem0210;
reg [WORD_WIDETH-1:0]           mem0211;
reg [WORD_WIDETH-1:0]           mem0212;
reg [WORD_WIDETH-1:0]           mem0213;
reg [WORD_WIDETH-1:0]           mem0214;
reg [WORD_WIDETH-1:0]           mem0215;
reg [WORD_WIDETH-1:0]           mem0216;
reg [WORD_WIDETH-1:0]           mem0217;
reg [WORD_WIDETH-1:0]           mem0218;
reg [WORD_WIDETH-1:0]           mem0300;
reg [WORD_WIDETH-1:0]           mem0301;
reg [WORD_WIDETH-1:0]           mem0302;
reg [WORD_WIDETH-1:0]           mem0303;
reg [WORD_WIDETH-1:0]           mem0304;
reg [WORD_WIDETH-1:0]           mem0305;
reg [WORD_WIDETH-1:0]           mem0306;
reg [WORD_WIDETH-1:0]           mem0307;
reg [WORD_WIDETH-1:0]           mem0308;
reg [WORD_WIDETH-1:0]           mem0309;
reg [WORD_WIDETH-1:0]           mem0310;
reg [WORD_WIDETH-1:0]           mem0311;
reg [WORD_WIDETH-1:0]           mem0312;
reg [WORD_WIDETH-1:0]           mem0313;
reg [WORD_WIDETH-1:0]           mem0314;
reg [WORD_WIDETH-1:0]           mem0315;
reg [WORD_WIDETH-1:0]           mem0316;
reg [WORD_WIDETH-1:0]           mem0317;
reg [WORD_WIDETH-1:0]           mem0318;
reg [WORD_WIDETH-1:0]           mem0400;
reg [WORD_WIDETH-1:0]           mem0401;
reg [WORD_WIDETH-1:0]           mem0402;
reg [WORD_WIDETH-1:0]           mem0403;
reg [WORD_WIDETH-1:0]           mem0404;
reg [WORD_WIDETH-1:0]           mem0405;
reg [WORD_WIDETH-1:0]           mem0406;
reg [WORD_WIDETH-1:0]           mem0407;
reg [WORD_WIDETH-1:0]           mem0408;
reg [WORD_WIDETH-1:0]           mem0409;
reg [WORD_WIDETH-1:0]           mem0410;
reg [WORD_WIDETH-1:0]           mem0411;
reg [WORD_WIDETH-1:0]           mem0412;
reg [WORD_WIDETH-1:0]           mem0413;
reg [WORD_WIDETH-1:0]           mem0414;
reg [WORD_WIDETH-1:0]           mem0415;
reg [WORD_WIDETH-1:0]           mem0416;
reg [WORD_WIDETH-1:0]           mem0417;
reg [WORD_WIDETH-1:0]           mem0418;
reg [WORD_WIDETH-1:0]           mem0500;
reg [WORD_WIDETH-1:0]           mem0501;
reg [WORD_WIDETH-1:0]           mem0502;
reg [WORD_WIDETH-1:0]           mem0503;
reg [WORD_WIDETH-1:0]           mem0504;
reg [WORD_WIDETH-1:0]           mem0505;
reg [WORD_WIDETH-1:0]           mem0506;
reg [WORD_WIDETH-1:0]           mem0507;
reg [WORD_WIDETH-1:0]           mem0508;
reg [WORD_WIDETH-1:0]           mem0509;
reg [WORD_WIDETH-1:0]           mem0510;
reg [WORD_WIDETH-1:0]           mem0511;
reg [WORD_WIDETH-1:0]           mem0512;
reg [WORD_WIDETH-1:0]           mem0513;
reg [WORD_WIDETH-1:0]           mem0514;
reg [WORD_WIDETH-1:0]           mem0515;
reg [WORD_WIDETH-1:0]           mem0516;
reg [WORD_WIDETH-1:0]           mem0517;
reg [WORD_WIDETH-1:0]           mem0518;
reg [WORD_WIDETH-1:0]           mem0600;
reg [WORD_WIDETH-1:0]           mem0601;
reg [WORD_WIDETH-1:0]           mem0602;
reg [WORD_WIDETH-1:0]           mem0603;
reg [WORD_WIDETH-1:0]           mem0604;
reg [WORD_WIDETH-1:0]           mem0605;
reg [WORD_WIDETH-1:0]           mem0606;
reg [WORD_WIDETH-1:0]           mem0607;
reg [WORD_WIDETH-1:0]           mem0608;
reg [WORD_WIDETH-1:0]           mem0609;
reg [WORD_WIDETH-1:0]           mem0610;
reg [WORD_WIDETH-1:0]           mem0611;
reg [WORD_WIDETH-1:0]           mem0612;
reg [WORD_WIDETH-1:0]           mem0613;
reg [WORD_WIDETH-1:0]           mem0614;
reg [WORD_WIDETH-1:0]           mem0615;
reg [WORD_WIDETH-1:0]           mem0616;
reg [WORD_WIDETH-1:0]           mem0617;
reg [WORD_WIDETH-1:0]           mem0618;
reg [WORD_WIDETH-1:0]           mem0700;
reg [WORD_WIDETH-1:0]           mem0701;
reg [WORD_WIDETH-1:0]           mem0702;
reg [WORD_WIDETH-1:0]           mem0703;
reg [WORD_WIDETH-1:0]           mem0704;
reg [WORD_WIDETH-1:0]           mem0705;
reg [WORD_WIDETH-1:0]           mem0706;
reg [WORD_WIDETH-1:0]           mem0707;
reg [WORD_WIDETH-1:0]           mem0708;
reg [WORD_WIDETH-1:0]           mem0709;
reg [WORD_WIDETH-1:0]           mem0710;
reg [WORD_WIDETH-1:0]           mem0711;
reg [WORD_WIDETH-1:0]           mem0712;
reg [WORD_WIDETH-1:0]           mem0713;
reg [WORD_WIDETH-1:0]           mem0714;
reg [WORD_WIDETH-1:0]           mem0715;
reg [WORD_WIDETH-1:0]           mem0716;
reg [WORD_WIDETH-1:0]           mem0717;
reg [WORD_WIDETH-1:0]           mem0718;
reg [WORD_WIDETH-1:0]           mem0800;
reg [WORD_WIDETH-1:0]           mem0801;
reg [WORD_WIDETH-1:0]           mem0802;
reg [WORD_WIDETH-1:0]           mem0803;
reg [WORD_WIDETH-1:0]           mem0804;
reg [WORD_WIDETH-1:0]           mem0805;
reg [WORD_WIDETH-1:0]           mem0806;
reg [WORD_WIDETH-1:0]           mem0807;
reg [WORD_WIDETH-1:0]           mem0808;
reg [WORD_WIDETH-1:0]           mem0809;
reg [WORD_WIDETH-1:0]           mem0810;
reg [WORD_WIDETH-1:0]           mem0811;
reg [WORD_WIDETH-1:0]           mem0812;
reg [WORD_WIDETH-1:0]           mem0813;
reg [WORD_WIDETH-1:0]           mem0814;
reg [WORD_WIDETH-1:0]           mem0815;
reg [WORD_WIDETH-1:0]           mem0816;
reg [WORD_WIDETH-1:0]           mem0817;
reg [WORD_WIDETH-1:0]           mem0818;
reg [WORD_WIDETH-1:0]           mem0900;
reg [WORD_WIDETH-1:0]           mem0901;
reg [WORD_WIDETH-1:0]           mem0902;
reg [WORD_WIDETH-1:0]           mem0903;
reg [WORD_WIDETH-1:0]           mem0904;
reg [WORD_WIDETH-1:0]           mem0905;
reg [WORD_WIDETH-1:0]           mem0906;
reg [WORD_WIDETH-1:0]           mem0907;
reg [WORD_WIDETH-1:0]           mem0908;
reg [WORD_WIDETH-1:0]           mem0909;
reg [WORD_WIDETH-1:0]           mem0910;
reg [WORD_WIDETH-1:0]           mem0911;
reg [WORD_WIDETH-1:0]           mem0912;
reg [WORD_WIDETH-1:0]           mem0913;
reg [WORD_WIDETH-1:0]           mem0914;
reg [WORD_WIDETH-1:0]           mem0915;
reg [WORD_WIDETH-1:0]           mem0916;
reg [WORD_WIDETH-1:0]           mem0917;
reg [WORD_WIDETH-1:0]           mem0918;
reg [WORD_WIDETH-1:0]           mem1000;
reg [WORD_WIDETH-1:0]           mem1001;
reg [WORD_WIDETH-1:0]           mem1002;
reg [WORD_WIDETH-1:0]           mem1003;
reg [WORD_WIDETH-1:0]           mem1004;
reg [WORD_WIDETH-1:0]           mem1005;
reg [WORD_WIDETH-1:0]           mem1006;
reg [WORD_WIDETH-1:0]           mem1007;
reg [WORD_WIDETH-1:0]           mem1008;
reg [WORD_WIDETH-1:0]           mem1009;
reg [WORD_WIDETH-1:0]           mem1010;
reg [WORD_WIDETH-1:0]           mem1011;
reg [WORD_WIDETH-1:0]           mem1012;
reg [WORD_WIDETH-1:0]           mem1013;
reg [WORD_WIDETH-1:0]           mem1014;
reg [WORD_WIDETH-1:0]           mem1015;
reg [WORD_WIDETH-1:0]           mem1016;
reg [WORD_WIDETH-1:0]           mem1017;
reg [WORD_WIDETH-1:0]           mem1018;
reg [WORD_WIDETH-1:0]           mem1100;
reg [WORD_WIDETH-1:0]           mem1101;
reg [WORD_WIDETH-1:0]           mem1102;
reg [WORD_WIDETH-1:0]           mem1103;
reg [WORD_WIDETH-1:0]           mem1104;
reg [WORD_WIDETH-1:0]           mem1105;
reg [WORD_WIDETH-1:0]           mem1106;
reg [WORD_WIDETH-1:0]           mem1107;
reg [WORD_WIDETH-1:0]           mem1108;
reg [WORD_WIDETH-1:0]           mem1109;
reg [WORD_WIDETH-1:0]           mem1110;
reg [WORD_WIDETH-1:0]           mem1111;
reg [WORD_WIDETH-1:0]           mem1112;
reg [WORD_WIDETH-1:0]           mem1113;
reg [WORD_WIDETH-1:0]           mem1114;
reg [WORD_WIDETH-1:0]           mem1115;
reg [WORD_WIDETH-1:0]           mem1116;
reg [WORD_WIDETH-1:0]           mem1117;
reg [WORD_WIDETH-1:0]           mem1118;
reg [WORD_WIDETH-1:0]           mem1200;
reg [WORD_WIDETH-1:0]           mem1201;
reg [WORD_WIDETH-1:0]           mem1202;
reg [WORD_WIDETH-1:0]           mem1203;
reg [WORD_WIDETH-1:0]           mem1204;
reg [WORD_WIDETH-1:0]           mem1205;
reg [WORD_WIDETH-1:0]           mem1206;
reg [WORD_WIDETH-1:0]           mem1207;
reg [WORD_WIDETH-1:0]           mem1208;
reg [WORD_WIDETH-1:0]           mem1209;
reg [WORD_WIDETH-1:0]           mem1210;
reg [WORD_WIDETH-1:0]           mem1211;
reg [WORD_WIDETH-1:0]           mem1212;
reg [WORD_WIDETH-1:0]           mem1213;
reg [WORD_WIDETH-1:0]           mem1214;
reg [WORD_WIDETH-1:0]           mem1215;
reg [WORD_WIDETH-1:0]           mem1216;
reg [WORD_WIDETH-1:0]           mem1217;
reg [WORD_WIDETH-1:0]           mem1218;
reg [WORD_WIDETH-1:0]           mem1300;
reg [WORD_WIDETH-1:0]           mem1301;
reg [WORD_WIDETH-1:0]           mem1302;
reg [WORD_WIDETH-1:0]           mem1303;
reg [WORD_WIDETH-1:0]           mem1304;
reg [WORD_WIDETH-1:0]           mem1305;
reg [WORD_WIDETH-1:0]           mem1306;
reg [WORD_WIDETH-1:0]           mem1307;
reg [WORD_WIDETH-1:0]           mem1308;
reg [WORD_WIDETH-1:0]           mem1309;
reg [WORD_WIDETH-1:0]           mem1310;
reg [WORD_WIDETH-1:0]           mem1311;
reg [WORD_WIDETH-1:0]           mem1312;
reg [WORD_WIDETH-1:0]           mem1313;
reg [WORD_WIDETH-1:0]           mem1314;
reg [WORD_WIDETH-1:0]           mem1315;
reg [WORD_WIDETH-1:0]           mem1316;
reg [WORD_WIDETH-1:0]           mem1317;
reg [WORD_WIDETH-1:0]           mem1318;
reg [WORD_WIDETH-1:0]           mem1400;
reg [WORD_WIDETH-1:0]           mem1401;
reg [WORD_WIDETH-1:0]           mem1402;
reg [WORD_WIDETH-1:0]           mem1403;
reg [WORD_WIDETH-1:0]           mem1404;
reg [WORD_WIDETH-1:0]           mem1405;
reg [WORD_WIDETH-1:0]           mem1406;
reg [WORD_WIDETH-1:0]           mem1407;
reg [WORD_WIDETH-1:0]           mem1408;
reg [WORD_WIDETH-1:0]           mem1409;
reg [WORD_WIDETH-1:0]           mem1410;
reg [WORD_WIDETH-1:0]           mem1411;
reg [WORD_WIDETH-1:0]           mem1412;
reg [WORD_WIDETH-1:0]           mem1413;
reg [WORD_WIDETH-1:0]           mem1414;
reg [WORD_WIDETH-1:0]           mem1415;
reg [WORD_WIDETH-1:0]           mem1416;
reg [WORD_WIDETH-1:0]           mem1417;
reg [WORD_WIDETH-1:0]           mem1418;
reg [WORD_WIDETH-1:0]           mem1500;
reg [WORD_WIDETH-1:0]           mem1501;
reg [WORD_WIDETH-1:0]           mem1502;
reg [WORD_WIDETH-1:0]           mem1503;
reg [WORD_WIDETH-1:0]           mem1504;
reg [WORD_WIDETH-1:0]           mem1505;
reg [WORD_WIDETH-1:0]           mem1506;
reg [WORD_WIDETH-1:0]           mem1507;
reg [WORD_WIDETH-1:0]           mem1508;
reg [WORD_WIDETH-1:0]           mem1509;
reg [WORD_WIDETH-1:0]           mem1510;
reg [WORD_WIDETH-1:0]           mem1511;
reg [WORD_WIDETH-1:0]           mem1512;
reg [WORD_WIDETH-1:0]           mem1513;
reg [WORD_WIDETH-1:0]           mem1514;
reg [WORD_WIDETH-1:0]           mem1515;
reg [WORD_WIDETH-1:0]           mem1516;
reg [WORD_WIDETH-1:0]           mem1517;
reg [WORD_WIDETH-1:0]           mem1518;
reg [WORD_WIDETH-1:0]           mem1600;
reg [WORD_WIDETH-1:0]           mem1601;
reg [WORD_WIDETH-1:0]           mem1602;
reg [WORD_WIDETH-1:0]           mem1603;
reg [WORD_WIDETH-1:0]           mem1604;
reg [WORD_WIDETH-1:0]           mem1605;
reg [WORD_WIDETH-1:0]           mem1606;
reg [WORD_WIDETH-1:0]           mem1607;
reg [WORD_WIDETH-1:0]           mem1608;
reg [WORD_WIDETH-1:0]           mem1609;
reg [WORD_WIDETH-1:0]           mem1610;
reg [WORD_WIDETH-1:0]           mem1611;
reg [WORD_WIDETH-1:0]           mem1612;
reg [WORD_WIDETH-1:0]           mem1613;
reg [WORD_WIDETH-1:0]           mem1614;
reg [WORD_WIDETH-1:0]           mem1615;
reg [WORD_WIDETH-1:0]           mem1616;
reg [WORD_WIDETH-1:0]           mem1617;
reg [WORD_WIDETH-1:0]           mem1618;
reg [WORD_WIDETH-1:0]           mem1700;
reg [WORD_WIDETH-1:0]           mem1701;
reg [WORD_WIDETH-1:0]           mem1702;
reg [WORD_WIDETH-1:0]           mem1703;
reg [WORD_WIDETH-1:0]           mem1704;
reg [WORD_WIDETH-1:0]           mem1705;
reg [WORD_WIDETH-1:0]           mem1706;
reg [WORD_WIDETH-1:0]           mem1707;
reg [WORD_WIDETH-1:0]           mem1708;
reg [WORD_WIDETH-1:0]           mem1709;
reg [WORD_WIDETH-1:0]           mem1710;
reg [WORD_WIDETH-1:0]           mem1711;
reg [WORD_WIDETH-1:0]           mem1712;
reg [WORD_WIDETH-1:0]           mem1713;
reg [WORD_WIDETH-1:0]           mem1714;
reg [WORD_WIDETH-1:0]           mem1715;
reg [WORD_WIDETH-1:0]           mem1716;
reg [WORD_WIDETH-1:0]           mem1717;
reg [WORD_WIDETH-1:0]           mem1718;
reg [WORD_WIDETH-1:0]           mem1800;
reg [WORD_WIDETH-1:0]           mem1801;
reg [WORD_WIDETH-1:0]           mem1802;
reg [WORD_WIDETH-1:0]           mem1803;
reg [WORD_WIDETH-1:0]           mem1804;
reg [WORD_WIDETH-1:0]           mem1805;
reg [WORD_WIDETH-1:0]           mem1806;
reg [WORD_WIDETH-1:0]           mem1807;
reg [WORD_WIDETH-1:0]           mem1808;
reg [WORD_WIDETH-1:0]           mem1809;
reg [WORD_WIDETH-1:0]           mem1810;
reg [WORD_WIDETH-1:0]           mem1811;
reg [WORD_WIDETH-1:0]           mem1812;
reg [WORD_WIDETH-1:0]           mem1813;
reg [WORD_WIDETH-1:0]           mem1814;
reg [WORD_WIDETH-1:0]           mem1815;
reg [WORD_WIDETH-1:0]           mem1816;
reg [WORD_WIDETH-1:0]           mem1817;
reg [WORD_WIDETH-1:0]           mem1818;

/**********************************************************************************************************************/
/************************INPUT Logic *********************************************************************************/
/**********************************************************************************************************************/
reg [WORD_WIDETH*19-1:0] input_buffer;
reg [23:0] input_extra_buffer;


/************************INPUT Logic END****************************/

/**********************************************************************************************************************/
/************************SWITCH Logic *********************************************************************************/
/**********************************************************************************************************************/
always @ (clk)
begin
    if(ctr_word==4'h1)
    begin
        mem0000 <= mem0400;
        mem0001 <= mem0401;
        mem0002 <= mem0402;
        mem0003 <= mem0403;
        mem0004 <= mem0404;
        mem0005 <= mem0405;
        mem0006 <= mem0406;
        mem0007 <= mem0407;
        mem0008 <= mem0408;
        mem0009 <= mem0409;
        mem0010 <= mem0410;
        mem0011 <= mem0411;
        mem0012 <= mem0412;
        mem0013 <= mem0413;
        mem0014 <= mem0414;
        mem0015 <= mem0415;
        mem0016 <= mem0416;
        mem0017 <= mem0417;
        mem0018 <= mem0418;
    end
    else
    begin
        mem0000 <= mem0000;
        mem0001 <= mem0001;
        mem0002 <= mem0002;
        mem0003 <= mem0003;
        mem0004 <= mem0004;
        mem0005 <= mem0005;
        mem0006 <= mem0006;
        mem0007 <= mem0007;
        mem0008 <= mem0008;
        mem0009 <= mem0009;
        mem0010 <= mem0010;
        mem0011 <= mem0011;
        mem0012 <= mem0012;
        mem0013 <= mem0013;
        mem0014 <= mem0014;
        mem0015 <= mem0015;
        mem0016 <= mem0016;
        mem0017 <= mem0017;
        mem0018 <= mem0018;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h2)
    begin
        mem0100 <= mem0500;
        mem0101 <= mem0501;
        mem0102 <= mem0502;
        mem0103 <= mem0503;
        mem0104 <= mem0504;
        mem0105 <= mem0505;
        mem0106 <= mem0506;
        mem0107 <= mem0507;
        mem0108 <= mem0508;
        mem0109 <= mem0509;
        mem0110 <= mem0510;
        mem0111 <= mem0511;
        mem0112 <= mem0512;
        mem0113 <= mem0513;
        mem0114 <= mem0514;
        mem0115 <= mem0515;
        mem0116 <= mem0516;
        mem0117 <= mem0517;
        mem0118 <= mem0518;
    end
    else
    begin
        mem0100 <= mem0100;
        mem0101 <= mem0101;
        mem0102 <= mem0102;
        mem0103 <= mem0103;
        mem0104 <= mem0104;
        mem0105 <= mem0105;
        mem0106 <= mem0106;
        mem0107 <= mem0107;
        mem0108 <= mem0108;
        mem0109 <= mem0109;
        mem0110 <= mem0110;
        mem0111 <= mem0111;
        mem0112 <= mem0112;
        mem0113 <= mem0113;
        mem0114 <= mem0114;
        mem0115 <= mem0115;
        mem0116 <= mem0116;
        mem0117 <= mem0117;
        mem0118 <= mem0118;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h3)
    begin
        mem0200 <= mem0600;
        mem0201 <= mem0601;
        mem0202 <= mem0602;
        mem0203 <= mem0603;
        mem0204 <= mem0604;
        mem0205 <= mem0605;
        mem0206 <= mem0606;
        mem0207 <= mem0607;
        mem0208 <= mem0608;
        mem0209 <= mem0609;
        mem0210 <= mem0610;
        mem0211 <= mem0611;
        mem0212 <= mem0612;
        mem0213 <= mem0613;
        mem0214 <= mem0614;
        mem0215 <= mem0615;
        mem0216 <= mem0616;
        mem0217 <= mem0617;
        mem0218 <= mem0618;
    end
    else
    begin
        mem0200 <= mem0200;
        mem0201 <= mem0201;
        mem0202 <= mem0202;
        mem0203 <= mem0203;
        mem0204 <= mem0204;
        mem0205 <= mem0205;
        mem0206 <= mem0206;
        mem0207 <= mem0207;
        mem0208 <= mem0208;
        mem0209 <= mem0209;
        mem0210 <= mem0210;
        mem0211 <= mem0211;
        mem0212 <= mem0212;
        mem0213 <= mem0213;
        mem0214 <= mem0214;
        mem0215 <= mem0215;
        mem0216 <= mem0216;
        mem0217 <= mem0217;
        mem0218 <= mem0218;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h4)
    begin
        mem0300 <= mem0700;
        mem0301 <= mem0701;
        mem0302 <= mem0702;
        mem0303 <= mem0703;
        mem0304 <= mem0704;
        mem0305 <= mem0705;
        mem0306 <= mem0706;
        mem0307 <= mem0707;
        mem0308 <= mem0708;
        mem0309 <= mem0709;
        mem0310 <= mem0710;
        mem0311 <= mem0711;
        mem0312 <= mem0712;
        mem0313 <= mem0713;
        mem0314 <= mem0714;
        mem0315 <= mem0715;
        mem0316 <= mem0716;
        mem0317 <= mem0717;
        mem0318 <= mem0718;
    end
    else
    begin
        mem0300 <= mem0300;
        mem0301 <= mem0301;
        mem0302 <= mem0302;
        mem0303 <= mem0303;
        mem0304 <= mem0304;
        mem0305 <= mem0305;
        mem0306 <= mem0306;
        mem0307 <= mem0307;
        mem0308 <= mem0308;
        mem0309 <= mem0309;
        mem0310 <= mem0310;
        mem0311 <= mem0311;
        mem0312 <= mem0312;
        mem0313 <= mem0313;
        mem0314 <= mem0314;
        mem0315 <= mem0315;
        mem0316 <= mem0316;
        mem0317 <= mem0317;
        mem0318 <= mem0318;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h5)
    begin
        mem0400 <= mem0800;
        mem0401 <= mem0801;
        mem0402 <= mem0802;
        mem0403 <= mem0803;
        mem0404 <= mem0804;
        mem0405 <= mem0805;
        mem0406 <= mem0806;
        mem0407 <= mem0807;
        mem0408 <= mem0808;
        mem0409 <= mem0809;
        mem0410 <= mem0810;
        mem0411 <= mem0811;
        mem0412 <= mem0812;
        mem0413 <= mem0813;
        mem0414 <= mem0814;
        mem0415 <= mem0815;
        mem0416 <= mem0816;
        mem0417 <= mem0817;
        mem0418 <= mem0818;
    end
    else
    begin
        mem0400 <= mem0400;
        mem0401 <= mem0401;
        mem0402 <= mem0402;
        mem0403 <= mem0403;
        mem0404 <= mem0404;
        mem0405 <= mem0405;
        mem0406 <= mem0406;
        mem0407 <= mem0407;
        mem0408 <= mem0408;
        mem0409 <= mem0409;
        mem0410 <= mem0410;
        mem0411 <= mem0411;
        mem0412 <= mem0412;
        mem0413 <= mem0413;
        mem0414 <= mem0414;
        mem0415 <= mem0415;
        mem0416 <= mem0416;
        mem0417 <= mem0417;
        mem0418 <= mem0418;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h6)
    begin
        mem0500 <= mem0900;
        mem0501 <= mem0901;
        mem0502 <= mem0902;
        mem0503 <= mem0903;
        mem0504 <= mem0904;
        mem0505 <= mem0905;
        mem0506 <= mem0906;
        mem0507 <= mem0907;
        mem0508 <= mem0908;
        mem0509 <= mem0909;
        mem0510 <= mem0910;
        mem0511 <= mem0911;
        mem0512 <= mem0912;
        mem0513 <= mem0913;
        mem0514 <= mem0914;
        mem0515 <= mem0915;
        mem0516 <= mem0916;
        mem0517 <= mem0917;
        mem0518 <= mem0918;
    end
    else
    begin
        mem0500 <= mem0500;
        mem0501 <= mem0501;
        mem0502 <= mem0502;
        mem0503 <= mem0503;
        mem0504 <= mem0504;
        mem0505 <= mem0505;
        mem0506 <= mem0506;
        mem0507 <= mem0507;
        mem0508 <= mem0508;
        mem0509 <= mem0509;
        mem0510 <= mem0510;
        mem0511 <= mem0511;
        mem0512 <= mem0512;
        mem0513 <= mem0513;
        mem0514 <= mem0514;
        mem0515 <= mem0515;
        mem0516 <= mem0516;
        mem0517 <= mem0517;
        mem0518 <= mem0518;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h7)
    begin
        mem0600 <= mem1000;
        mem0601 <= mem1001;
        mem0602 <= mem1002;
        mem0603 <= mem1003;
        mem0604 <= mem1004;
        mem0605 <= mem1005;
        mem0606 <= mem1006;
        mem0607 <= mem1007;
        mem0608 <= mem1008;
        mem0609 <= mem1009;
        mem0610 <= mem1010;
        mem0611 <= mem1011;
        mem0612 <= mem1012;
        mem0613 <= mem1013;
        mem0614 <= mem1014;
        mem0615 <= mem1015;
        mem0616 <= mem1016;
        mem0617 <= mem1017;
        mem0618 <= mem1018;
    end
    else
    begin
        mem0600 <= mem0600;
        mem0601 <= mem0601;
        mem0602 <= mem0602;
        mem0603 <= mem0603;
        mem0604 <= mem0604;
        mem0605 <= mem0605;
        mem0606 <= mem0606;
        mem0607 <= mem0607;
        mem0608 <= mem0608;
        mem0609 <= mem0609;
        mem0610 <= mem0610;
        mem0611 <= mem0611;
        mem0612 <= mem0612;
        mem0613 <= mem0613;
        mem0614 <= mem0614;
        mem0615 <= mem0615;
        mem0616 <= mem0616;
        mem0617 <= mem0617;
        mem0618 <= mem0618;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h8)
    begin
        mem0700 <= mem1100;
        mem0701 <= mem1101;
        mem0702 <= mem1102;
        mem0703 <= mem1103;
        mem0704 <= mem1104;
        mem0705 <= mem1105;
        mem0706 <= mem1106;
        mem0707 <= mem1107;
        mem0708 <= mem1108;
        mem0709 <= mem1109;
        mem0710 <= mem1110;
        mem0711 <= mem1111;
        mem0712 <= mem1112;
        mem0713 <= mem1113;
        mem0714 <= mem1114;
        mem0715 <= mem1115;
        mem0716 <= mem1116;
        mem0717 <= mem1117;
        mem0718 <= mem1118;
    end
    else
    begin
        mem0700 <= mem0700;
        mem0701 <= mem0701;
        mem0702 <= mem0702;
        mem0703 <= mem0703;
        mem0704 <= mem0704;
        mem0705 <= mem0705;
        mem0706 <= mem0706;
        mem0707 <= mem0707;
        mem0708 <= mem0708;
        mem0709 <= mem0709;
        mem0710 <= mem0710;
        mem0711 <= mem0711;
        mem0712 <= mem0712;
        mem0713 <= mem0713;
        mem0714 <= mem0714;
        mem0715 <= mem0715;
        mem0716 <= mem0716;
        mem0717 <= mem0717;
        mem0718 <= mem0718;
    end
end

always @ (clk)
begin
    if(ctr_word==4'h9)
    begin
        mem0800 <= mem1200;
        mem0801 <= mem1201;
        mem0802 <= mem1202;
        mem0803 <= mem1203;
        mem0804 <= mem1204;
        mem0805 <= mem1205;
        mem0806 <= mem1206;
        mem0807 <= mem1207;
        mem0808 <= mem1208;
        mem0809 <= mem1209;
        mem0810 <= mem1210;
        mem0811 <= mem1211;
        mem0812 <= mem1212;
        mem0813 <= mem1213;
        mem0814 <= mem1214;
        mem0815 <= mem1215;
        mem0816 <= mem1216;
        mem0817 <= mem1217;
        mem0818 <= mem1218;
    end
    else
    begin
        mem0800 <= mem0800;
        mem0801 <= mem0801;
        mem0802 <= mem0802;
        mem0803 <= mem0803;
        mem0804 <= mem0804;
        mem0805 <= mem0805;
        mem0806 <= mem0806;
        mem0807 <= mem0807;
        mem0808 <= mem0808;
        mem0809 <= mem0809;
        mem0810 <= mem0810;
        mem0811 <= mem0811;
        mem0812 <= mem0812;
        mem0813 <= mem0813;
        mem0814 <= mem0814;
        mem0815 <= mem0815;
        mem0816 <= mem0816;
        mem0817 <= mem0817;
        mem0818 <= mem0818;
    end
end

always @ (clk)
begin
    if(ctr_word==4'ha)
    begin
        mem0900 <= mem1300;
        mem0901 <= mem1301;
        mem0902 <= mem1302;
        mem0903 <= mem1303;
        mem0904 <= mem1304;
        mem0905 <= mem1305;
        mem0906 <= mem1306;
        mem0907 <= mem1307;
        mem0908 <= mem1308;
        mem0909 <= mem1309;
        mem0910 <= mem1310;
        mem0911 <= mem1311;
        mem0912 <= mem1312;
        mem0913 <= mem1313;
        mem0914 <= mem1314;
        mem0915 <= mem1315;
        mem0916 <= mem1316;
        mem0917 <= mem1317;
        mem0918 <= mem1318;
    end
    else
    begin
        mem0900 <= mem0900;
        mem0901 <= mem0901;
        mem0902 <= mem0902;
        mem0903 <= mem0903;
        mem0904 <= mem0904;
        mem0905 <= mem0905;
        mem0906 <= mem0906;
        mem0907 <= mem0907;
        mem0908 <= mem0908;
        mem0909 <= mem0909;
        mem0910 <= mem0910;
        mem0911 <= mem0911;
        mem0912 <= mem0912;
        mem0913 <= mem0913;
        mem0914 <= mem0914;
        mem0915 <= mem0915;
        mem0916 <= mem0916;
        mem0917 <= mem0917;
        mem0918 <= mem0918;
    end
end

always @ (clk)
begin
    if(ctr_word==4'hb)
    begin
        mem1000 <= mem1400;
        mem1001 <= mem1401;
        mem1002 <= mem1402;
        mem1003 <= mem1403;
        mem1004 <= mem1404;
        mem1005 <= mem1405;
        mem1006 <= mem1406;
        mem1007 <= mem1407;
        mem1008 <= mem1408;
        mem1009 <= mem1409;
        mem1010 <= mem1410;
        mem1011 <= mem1411;
        mem1012 <= mem1412;
        mem1013 <= mem1413;
        mem1014 <= mem1414;
        mem1015 <= mem1415;
        mem1016 <= mem1416;
        mem1017 <= mem1417;
        mem1018 <= mem1418;
    end
    else
    begin
        mem1000 <= mem1000;
        mem1001 <= mem1001;
        mem1002 <= mem1002;
        mem1003 <= mem1003;
        mem1004 <= mem1004;
        mem1005 <= mem1005;
        mem1006 <= mem1006;
        mem1007 <= mem1007;
        mem1008 <= mem1008;
        mem1009 <= mem1009;
        mem1010 <= mem1010;
        mem1011 <= mem1011;
        mem1012 <= mem1012;
        mem1013 <= mem1013;
        mem1014 <= mem1014;
        mem1015 <= mem1015;
        mem1016 <= mem1016;
        mem1017 <= mem1017;
        mem1018 <= mem1018;
    end
end

always @ (clk)
begin
    if(ctr_word==4'hc)
    begin
        mem1100 <= mem1500;
        mem1101 <= mem1501;
        mem1102 <= mem1502;
        mem1103 <= mem1503;
        mem1104 <= mem1504;
        mem1105 <= mem1505;
        mem1106 <= mem1506;
        mem1107 <= mem1507;
        mem1108 <= mem1508;
        mem1109 <= mem1509;
        mem1110 <= mem1510;
        mem1111 <= mem1511;
        mem1112 <= mem1512;
        mem1113 <= mem1513;
        mem1114 <= mem1514;
        mem1115 <= mem1515;
        mem1116 <= mem1516;
        mem1117 <= mem1517;
        mem1118 <= mem1518;
    end
    else
    begin
        mem1100 <= mem1100;
        mem1101 <= mem1101;
        mem1102 <= mem1102;
        mem1103 <= mem1103;
        mem1104 <= mem1104;
        mem1105 <= mem1105;
        mem1106 <= mem1106;
        mem1107 <= mem1107;
        mem1108 <= mem1108;
        mem1109 <= mem1109;
        mem1110 <= mem1110;
        mem1111 <= mem1111;
        mem1112 <= mem1112;
        mem1113 <= mem1113;
        mem1114 <= mem1114;
        mem1115 <= mem1115;
        mem1116 <= mem1116;
        mem1117 <= mem1117;
        mem1118 <= mem1118;
    end
end

always @ (clk)
begin
    if(ctr_word==4'hd)
    begin
        mem1200 <= mem1600;
        mem1201 <= mem1601;
        mem1202 <= mem1602;
        mem1203 <= mem1603;
        mem1204 <= mem1604;
        mem1205 <= mem1605;
        mem1206 <= mem1606;
        mem1207 <= mem1607;
        mem1208 <= mem1608;
        mem1209 <= mem1609;
        mem1210 <= mem1610;
        mem1211 <= mem1611;
        mem1212 <= mem1612;
        mem1213 <= mem1613;
        mem1214 <= mem1614;
        mem1215 <= mem1615;
        mem1216 <= mem1616;
        mem1217 <= mem1617;
        mem1218 <= mem1618;
    end
    else
    begin
        mem1200 <= mem1200;
        mem1201 <= mem1201;
        mem1202 <= mem1202;
        mem1203 <= mem1203;
        mem1204 <= mem1204;
        mem1205 <= mem1205;
        mem1206 <= mem1206;
        mem1207 <= mem1207;
        mem1208 <= mem1208;
        mem1209 <= mem1209;
        mem1210 <= mem1210;
        mem1211 <= mem1211;
        mem1212 <= mem1212;
        mem1213 <= mem1213;
        mem1214 <= mem1214;
        mem1215 <= mem1215;
        mem1216 <= mem1216;
        mem1217 <= mem1217;
        mem1218 <= mem1218;
    end
end

always @ (clk)
begin
    if(ctr_word==4'he)
    begin
        mem1300 <= mem1700;
        mem1301 <= mem1701;
        mem1302 <= mem1702;
        mem1303 <= mem1703;
        mem1304 <= mem1704;
        mem1305 <= mem1705;
        mem1306 <= mem1706;
        mem1307 <= mem1707;
        mem1308 <= mem1708;
        mem1309 <= mem1709;
        mem1310 <= mem1710;
        mem1311 <= mem1711;
        mem1312 <= mem1712;
        mem1313 <= mem1713;
        mem1314 <= mem1714;
        mem1315 <= mem1715;
        mem1316 <= mem1716;
        mem1317 <= mem1717;
        mem1318 <= mem1718;
    end
    else
    begin
        mem1300 <= mem1300;
        mem1301 <= mem1301;
        mem1302 <= mem1302;
        mem1303 <= mem1303;
        mem1304 <= mem1304;
        mem1305 <= mem1305;
        mem1306 <= mem1306;
        mem1307 <= mem1307;
        mem1308 <= mem1308;
        mem1309 <= mem1309;
        mem1310 <= mem1310;
        mem1311 <= mem1311;
        mem1312 <= mem1312;
        mem1313 <= mem1313;
        mem1314 <= mem1314;
        mem1315 <= mem1315;
        mem1316 <= mem1316;
        mem1317 <= mem1317;
        mem1318 <= mem1318;
    end
end

always @ (clk)
begin
    if(ctr_word==4'hf)
    begin
        mem1400 <= mem1800;
        mem1401 <= mem1801;
        mem1402 <= mem1802;
        mem1403 <= mem1803;
        mem1404 <= mem1804;
        mem1405 <= mem1805;
        mem1406 <= mem1806;
        mem1407 <= mem1807;
        mem1408 <= mem1808;
        mem1409 <= mem1809;
        mem1410 <= mem1810;
        mem1411 <= mem1811;
        mem1412 <= mem1812;
        mem1413 <= mem1813;
        mem1414 <= mem1814;
        mem1415 <= mem1815;
        mem1416 <= mem1816;
        mem1417 <= mem1817;
        mem1418 <= mem1818;
    end
    else
    begin
        mem1400 <= mem1400;
        mem1401 <= mem1401;
        mem1402 <= mem1402;
        mem1403 <= mem1403;
        mem1404 <= mem1404;
        mem1405 <= mem1405;
        mem1406 <= mem1406;
        mem1407 <= mem1407;
        mem1408 <= mem1408;
        mem1409 <= mem1409;
        mem1410 <= mem1410;
        mem1411 <= mem1411;
        mem1412 <= mem1412;
        mem1413 <= mem1413;
        mem1414 <= mem1414;
        mem1415 <= mem1415;
        mem1416 <= mem1416;
        mem1417 <= mem1417;
        mem1418 <= mem1418;
    end
end


/************************SWITCH Logic END*******************/

/**********************************************************************************************************************/
/************************OUTPUT Logic *********************************************************************************/
/**********************************************************************************************************************/
always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in00 <= mem0000;
    4'h1: pe00_in00 <= mem0100;
    4'h2: pe00_in00 <= mem0200;
    4'h3: pe00_in00 <= mem0300;
    4'h4: pe00_in00 <= mem0400;
    4'h5: pe00_in00 <= mem0500;
    4'h6: pe00_in00 <= mem0600;
    4'h7: pe00_in00 <= mem0700;
    4'h8: pe00_in00 <= mem0800;
    4'h9: pe00_in00 <= mem0900;
    4'ha: pe00_in00 <= mem1000;
    4'hb: pe00_in00 <= mem1100;
    4'hc: pe00_in00 <= mem1200;
    4'hd: pe00_in00 <= mem1300;
    4'he: pe00_in00 <= mem1400;
    4'hf: pe00_in00 <= mem1500;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in01 <= mem0001;
    4'h1: pe00_in01 <= mem0101;
    4'h2: pe00_in01 <= mem0201;
    4'h3: pe00_in01 <= mem0301;
    4'h4: pe00_in01 <= mem0401;
    4'h5: pe00_in01 <= mem0501;
    4'h6: pe00_in01 <= mem0601;
    4'h7: pe00_in01 <= mem0701;
    4'h8: pe00_in01 <= mem0801;
    4'h9: pe00_in01 <= mem0901;
    4'ha: pe00_in01 <= mem1001;
    4'hb: pe00_in01 <= mem1101;
    4'hc: pe00_in01 <= mem1201;
    4'hd: pe00_in01 <= mem1301;
    4'he: pe00_in01 <= mem1401;
    4'hf: pe00_in01 <= mem1501;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in02 <= mem0002;
    4'h1: pe00_in02 <= mem0102;
    4'h2: pe00_in02 <= mem0202;
    4'h3: pe00_in02 <= mem0302;
    4'h4: pe00_in02 <= mem0402;
    4'h5: pe00_in02 <= mem0502;
    4'h6: pe00_in02 <= mem0602;
    4'h7: pe00_in02 <= mem0702;
    4'h8: pe00_in02 <= mem0802;
    4'h9: pe00_in02 <= mem0902;
    4'ha: pe00_in02 <= mem1002;
    4'hb: pe00_in02 <= mem1102;
    4'hc: pe00_in02 <= mem1202;
    4'hd: pe00_in02 <= mem1302;
    4'he: pe00_in02 <= mem1402;
    4'hf: pe00_in02 <= mem1502;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in03 <= mem0003;
    4'h1: pe00_in03 <= mem0103;
    4'h2: pe00_in03 <= mem0203;
    4'h3: pe00_in03 <= mem0303;
    4'h4: pe00_in03 <= mem0403;
    4'h5: pe00_in03 <= mem0503;
    4'h6: pe00_in03 <= mem0603;
    4'h7: pe00_in03 <= mem0703;
    4'h8: pe00_in03 <= mem0803;
    4'h9: pe00_in03 <= mem0903;
    4'ha: pe00_in03 <= mem1003;
    4'hb: pe00_in03 <= mem1103;
    4'hc: pe00_in03 <= mem1203;
    4'hd: pe00_in03 <= mem1303;
    4'he: pe00_in03 <= mem1403;
    4'hf: pe00_in03 <= mem1503;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in04 <= mem0100;
    4'h1: pe00_in04 <= mem0200;
    4'h2: pe00_in04 <= mem0300;
    4'h3: pe00_in04 <= mem0400;
    4'h4: pe00_in04 <= mem0500;
    4'h5: pe00_in04 <= mem0600;
    4'h6: pe00_in04 <= mem0700;
    4'h7: pe00_in04 <= mem0800;
    4'h8: pe00_in04 <= mem0900;
    4'h9: pe00_in04 <= mem1000;
    4'ha: pe00_in04 <= mem1100;
    4'hb: pe00_in04 <= mem1200;
    4'hc: pe00_in04 <= mem1300;
    4'hd: pe00_in04 <= mem1400;
    4'he: pe00_in04 <= mem1500;
    4'hf: pe00_in04 <= mem1600;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in05 <= mem0101;
    4'h1: pe00_in05 <= mem0201;
    4'h2: pe00_in05 <= mem0301;
    4'h3: pe00_in05 <= mem0401;
    4'h4: pe00_in05 <= mem0501;
    4'h5: pe00_in05 <= mem0601;
    4'h6: pe00_in05 <= mem0701;
    4'h7: pe00_in05 <= mem0801;
    4'h8: pe00_in05 <= mem0901;
    4'h9: pe00_in05 <= mem1001;
    4'ha: pe00_in05 <= mem1101;
    4'hb: pe00_in05 <= mem1201;
    4'hc: pe00_in05 <= mem1301;
    4'hd: pe00_in05 <= mem1401;
    4'he: pe00_in05 <= mem1501;
    4'hf: pe00_in05 <= mem1601;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in06 <= mem0102;
    4'h1: pe00_in06 <= mem0202;
    4'h2: pe00_in06 <= mem0302;
    4'h3: pe00_in06 <= mem0402;
    4'h4: pe00_in06 <= mem0502;
    4'h5: pe00_in06 <= mem0602;
    4'h6: pe00_in06 <= mem0702;
    4'h7: pe00_in06 <= mem0802;
    4'h8: pe00_in06 <= mem0902;
    4'h9: pe00_in06 <= mem1002;
    4'ha: pe00_in06 <= mem1102;
    4'hb: pe00_in06 <= mem1202;
    4'hc: pe00_in06 <= mem1302;
    4'hd: pe00_in06 <= mem1402;
    4'he: pe00_in06 <= mem1502;
    4'hf: pe00_in06 <= mem1602;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in07 <= mem0103;
    4'h1: pe00_in07 <= mem0203;
    4'h2: pe00_in07 <= mem0303;
    4'h3: pe00_in07 <= mem0403;
    4'h4: pe00_in07 <= mem0503;
    4'h5: pe00_in07 <= mem0603;
    4'h6: pe00_in07 <= mem0703;
    4'h7: pe00_in07 <= mem0803;
    4'h8: pe00_in07 <= mem0903;
    4'h9: pe00_in07 <= mem1003;
    4'ha: pe00_in07 <= mem1103;
    4'hb: pe00_in07 <= mem1203;
    4'hc: pe00_in07 <= mem1303;
    4'hd: pe00_in07 <= mem1403;
    4'he: pe00_in07 <= mem1503;
    4'hf: pe00_in07 <= mem1603;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in08 <= mem0200;
    4'h1: pe00_in08 <= mem0300;
    4'h2: pe00_in08 <= mem0400;
    4'h3: pe00_in08 <= mem0500;
    4'h4: pe00_in08 <= mem0600;
    4'h5: pe00_in08 <= mem0700;
    4'h6: pe00_in08 <= mem0800;
    4'h7: pe00_in08 <= mem0900;
    4'h8: pe00_in08 <= mem1000;
    4'h9: pe00_in08 <= mem1100;
    4'ha: pe00_in08 <= mem1200;
    4'hb: pe00_in08 <= mem1300;
    4'hc: pe00_in08 <= mem1400;
    4'hd: pe00_in08 <= mem1500;
    4'he: pe00_in08 <= mem1600;
    4'hf: pe00_in08 <= mem1700;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in09 <= mem0201;
    4'h1: pe00_in09 <= mem0301;
    4'h2: pe00_in09 <= mem0401;
    4'h3: pe00_in09 <= mem0501;
    4'h4: pe00_in09 <= mem0601;
    4'h5: pe00_in09 <= mem0701;
    4'h6: pe00_in09 <= mem0801;
    4'h7: pe00_in09 <= mem0901;
    4'h8: pe00_in09 <= mem1001;
    4'h9: pe00_in09 <= mem1101;
    4'ha: pe00_in09 <= mem1201;
    4'hb: pe00_in09 <= mem1301;
    4'hc: pe00_in09 <= mem1401;
    4'hd: pe00_in09 <= mem1501;
    4'he: pe00_in09 <= mem1601;
    4'hf: pe00_in09 <= mem1701;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in10 <= mem0202;
    4'h1: pe00_in10 <= mem0302;
    4'h2: pe00_in10 <= mem0402;
    4'h3: pe00_in10 <= mem0502;
    4'h4: pe00_in10 <= mem0602;
    4'h5: pe00_in10 <= mem0702;
    4'h6: pe00_in10 <= mem0802;
    4'h7: pe00_in10 <= mem0902;
    4'h8: pe00_in10 <= mem1002;
    4'h9: pe00_in10 <= mem1102;
    4'ha: pe00_in10 <= mem1202;
    4'hb: pe00_in10 <= mem1302;
    4'hc: pe00_in10 <= mem1402;
    4'hd: pe00_in10 <= mem1502;
    4'he: pe00_in10 <= mem1602;
    4'hf: pe00_in10 <= mem1702;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in11 <= mem0203;
    4'h1: pe00_in11 <= mem0303;
    4'h2: pe00_in11 <= mem0403;
    4'h3: pe00_in11 <= mem0503;
    4'h4: pe00_in11 <= mem0603;
    4'h5: pe00_in11 <= mem0703;
    4'h6: pe00_in11 <= mem0803;
    4'h7: pe00_in11 <= mem0903;
    4'h8: pe00_in11 <= mem1003;
    4'h9: pe00_in11 <= mem1103;
    4'ha: pe00_in11 <= mem1203;
    4'hb: pe00_in11 <= mem1303;
    4'hc: pe00_in11 <= mem1403;
    4'hd: pe00_in11 <= mem1503;
    4'he: pe00_in11 <= mem1603;
    4'hf: pe00_in11 <= mem1703;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in12 <= mem0300;
    4'h1: pe00_in12 <= mem0400;
    4'h2: pe00_in12 <= mem0500;
    4'h3: pe00_in12 <= mem0600;
    4'h4: pe00_in12 <= mem0700;
    4'h5: pe00_in12 <= mem0800;
    4'h6: pe00_in12 <= mem0900;
    4'h7: pe00_in12 <= mem1000;
    4'h8: pe00_in12 <= mem1100;
    4'h9: pe00_in12 <= mem1200;
    4'ha: pe00_in12 <= mem1300;
    4'hb: pe00_in12 <= mem1400;
    4'hc: pe00_in12 <= mem1500;
    4'hd: pe00_in12 <= mem1600;
    4'he: pe00_in12 <= mem1700;
    4'hf: pe00_in12 <= mem1800;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in13 <= mem0301;
    4'h1: pe00_in13 <= mem0401;
    4'h2: pe00_in13 <= mem0501;
    4'h3: pe00_in13 <= mem0601;
    4'h4: pe00_in13 <= mem0701;
    4'h5: pe00_in13 <= mem0801;
    4'h6: pe00_in13 <= mem0901;
    4'h7: pe00_in13 <= mem1001;
    4'h8: pe00_in13 <= mem1101;
    4'h9: pe00_in13 <= mem1201;
    4'ha: pe00_in13 <= mem1301;
    4'hb: pe00_in13 <= mem1401;
    4'hc: pe00_in13 <= mem1501;
    4'hd: pe00_in13 <= mem1601;
    4'he: pe00_in13 <= mem1701;
    4'hf: pe00_in13 <= mem1801;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in14 <= mem0302;
    4'h1: pe00_in14 <= mem0402;
    4'h2: pe00_in14 <= mem0502;
    4'h3: pe00_in14 <= mem0602;
    4'h4: pe00_in14 <= mem0702;
    4'h5: pe00_in14 <= mem0802;
    4'h6: pe00_in14 <= mem0902;
    4'h7: pe00_in14 <= mem1002;
    4'h8: pe00_in14 <= mem1102;
    4'h9: pe00_in14 <= mem1202;
    4'ha: pe00_in14 <= mem1302;
    4'hb: pe00_in14 <= mem1402;
    4'hc: pe00_in14 <= mem1502;
    4'hd: pe00_in14 <= mem1602;
    4'he: pe00_in14 <= mem1702;
    4'hf: pe00_in14 <= mem1802;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe00_in15 <= mem0303;
    4'h1: pe00_in15 <= mem0403;
    4'h2: pe00_in15 <= mem0503;
    4'h3: pe00_in15 <= mem0603;
    4'h4: pe00_in15 <= mem0703;
    4'h5: pe00_in15 <= mem0803;
    4'h6: pe00_in15 <= mem0903;
    4'h7: pe00_in15 <= mem1003;
    4'h8: pe00_in15 <= mem1103;
    4'h9: pe00_in15 <= mem1203;
    4'ha: pe00_in15 <= mem1303;
    4'hb: pe00_in15 <= mem1403;
    4'hc: pe00_in15 <= mem1503;
    4'hd: pe00_in15 <= mem1603;
    4'he: pe00_in15 <= mem1703;
    4'hf: pe00_in15 <= mem1803;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in00 <= mem0001;
    4'h1: pe01_in00 <= mem0101;
    4'h2: pe01_in00 <= mem0201;
    4'h3: pe01_in00 <= mem0301;
    4'h4: pe01_in00 <= mem0401;
    4'h5: pe01_in00 <= mem0501;
    4'h6: pe01_in00 <= mem0601;
    4'h7: pe01_in00 <= mem0701;
    4'h8: pe01_in00 <= mem0801;
    4'h9: pe01_in00 <= mem0901;
    4'ha: pe01_in00 <= mem1001;
    4'hb: pe01_in00 <= mem1101;
    4'hc: pe01_in00 <= mem1201;
    4'hd: pe01_in00 <= mem1301;
    4'he: pe01_in00 <= mem1401;
    4'hf: pe01_in00 <= mem1501;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in01 <= mem0002;
    4'h1: pe01_in01 <= mem0102;
    4'h2: pe01_in01 <= mem0202;
    4'h3: pe01_in01 <= mem0302;
    4'h4: pe01_in01 <= mem0402;
    4'h5: pe01_in01 <= mem0502;
    4'h6: pe01_in01 <= mem0602;
    4'h7: pe01_in01 <= mem0702;
    4'h8: pe01_in01 <= mem0802;
    4'h9: pe01_in01 <= mem0902;
    4'ha: pe01_in01 <= mem1002;
    4'hb: pe01_in01 <= mem1102;
    4'hc: pe01_in01 <= mem1202;
    4'hd: pe01_in01 <= mem1302;
    4'he: pe01_in01 <= mem1402;
    4'hf: pe01_in01 <= mem1502;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in02 <= mem0003;
    4'h1: pe01_in02 <= mem0103;
    4'h2: pe01_in02 <= mem0203;
    4'h3: pe01_in02 <= mem0303;
    4'h4: pe01_in02 <= mem0403;
    4'h5: pe01_in02 <= mem0503;
    4'h6: pe01_in02 <= mem0603;
    4'h7: pe01_in02 <= mem0703;
    4'h8: pe01_in02 <= mem0803;
    4'h9: pe01_in02 <= mem0903;
    4'ha: pe01_in02 <= mem1003;
    4'hb: pe01_in02 <= mem1103;
    4'hc: pe01_in02 <= mem1203;
    4'hd: pe01_in02 <= mem1303;
    4'he: pe01_in02 <= mem1403;
    4'hf: pe01_in02 <= mem1503;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in03 <= mem0004;
    4'h1: pe01_in03 <= mem0104;
    4'h2: pe01_in03 <= mem0204;
    4'h3: pe01_in03 <= mem0304;
    4'h4: pe01_in03 <= mem0404;
    4'h5: pe01_in03 <= mem0504;
    4'h6: pe01_in03 <= mem0604;
    4'h7: pe01_in03 <= mem0704;
    4'h8: pe01_in03 <= mem0804;
    4'h9: pe01_in03 <= mem0904;
    4'ha: pe01_in03 <= mem1004;
    4'hb: pe01_in03 <= mem1104;
    4'hc: pe01_in03 <= mem1204;
    4'hd: pe01_in03 <= mem1304;
    4'he: pe01_in03 <= mem1404;
    4'hf: pe01_in03 <= mem1504;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in04 <= mem0101;
    4'h1: pe01_in04 <= mem0201;
    4'h2: pe01_in04 <= mem0301;
    4'h3: pe01_in04 <= mem0401;
    4'h4: pe01_in04 <= mem0501;
    4'h5: pe01_in04 <= mem0601;
    4'h6: pe01_in04 <= mem0701;
    4'h7: pe01_in04 <= mem0801;
    4'h8: pe01_in04 <= mem0901;
    4'h9: pe01_in04 <= mem1001;
    4'ha: pe01_in04 <= mem1101;
    4'hb: pe01_in04 <= mem1201;
    4'hc: pe01_in04 <= mem1301;
    4'hd: pe01_in04 <= mem1401;
    4'he: pe01_in04 <= mem1501;
    4'hf: pe01_in04 <= mem1601;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in05 <= mem0102;
    4'h1: pe01_in05 <= mem0202;
    4'h2: pe01_in05 <= mem0302;
    4'h3: pe01_in05 <= mem0402;
    4'h4: pe01_in05 <= mem0502;
    4'h5: pe01_in05 <= mem0602;
    4'h6: pe01_in05 <= mem0702;
    4'h7: pe01_in05 <= mem0802;
    4'h8: pe01_in05 <= mem0902;
    4'h9: pe01_in05 <= mem1002;
    4'ha: pe01_in05 <= mem1102;
    4'hb: pe01_in05 <= mem1202;
    4'hc: pe01_in05 <= mem1302;
    4'hd: pe01_in05 <= mem1402;
    4'he: pe01_in05 <= mem1502;
    4'hf: pe01_in05 <= mem1602;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in06 <= mem0103;
    4'h1: pe01_in06 <= mem0203;
    4'h2: pe01_in06 <= mem0303;
    4'h3: pe01_in06 <= mem0403;
    4'h4: pe01_in06 <= mem0503;
    4'h5: pe01_in06 <= mem0603;
    4'h6: pe01_in06 <= mem0703;
    4'h7: pe01_in06 <= mem0803;
    4'h8: pe01_in06 <= mem0903;
    4'h9: pe01_in06 <= mem1003;
    4'ha: pe01_in06 <= mem1103;
    4'hb: pe01_in06 <= mem1203;
    4'hc: pe01_in06 <= mem1303;
    4'hd: pe01_in06 <= mem1403;
    4'he: pe01_in06 <= mem1503;
    4'hf: pe01_in06 <= mem1603;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in07 <= mem0104;
    4'h1: pe01_in07 <= mem0204;
    4'h2: pe01_in07 <= mem0304;
    4'h3: pe01_in07 <= mem0404;
    4'h4: pe01_in07 <= mem0504;
    4'h5: pe01_in07 <= mem0604;
    4'h6: pe01_in07 <= mem0704;
    4'h7: pe01_in07 <= mem0804;
    4'h8: pe01_in07 <= mem0904;
    4'h9: pe01_in07 <= mem1004;
    4'ha: pe01_in07 <= mem1104;
    4'hb: pe01_in07 <= mem1204;
    4'hc: pe01_in07 <= mem1304;
    4'hd: pe01_in07 <= mem1404;
    4'he: pe01_in07 <= mem1504;
    4'hf: pe01_in07 <= mem1604;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in08 <= mem0201;
    4'h1: pe01_in08 <= mem0301;
    4'h2: pe01_in08 <= mem0401;
    4'h3: pe01_in08 <= mem0501;
    4'h4: pe01_in08 <= mem0601;
    4'h5: pe01_in08 <= mem0701;
    4'h6: pe01_in08 <= mem0801;
    4'h7: pe01_in08 <= mem0901;
    4'h8: pe01_in08 <= mem1001;
    4'h9: pe01_in08 <= mem1101;
    4'ha: pe01_in08 <= mem1201;
    4'hb: pe01_in08 <= mem1301;
    4'hc: pe01_in08 <= mem1401;
    4'hd: pe01_in08 <= mem1501;
    4'he: pe01_in08 <= mem1601;
    4'hf: pe01_in08 <= mem1701;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in09 <= mem0202;
    4'h1: pe01_in09 <= mem0302;
    4'h2: pe01_in09 <= mem0402;
    4'h3: pe01_in09 <= mem0502;
    4'h4: pe01_in09 <= mem0602;
    4'h5: pe01_in09 <= mem0702;
    4'h6: pe01_in09 <= mem0802;
    4'h7: pe01_in09 <= mem0902;
    4'h8: pe01_in09 <= mem1002;
    4'h9: pe01_in09 <= mem1102;
    4'ha: pe01_in09 <= mem1202;
    4'hb: pe01_in09 <= mem1302;
    4'hc: pe01_in09 <= mem1402;
    4'hd: pe01_in09 <= mem1502;
    4'he: pe01_in09 <= mem1602;
    4'hf: pe01_in09 <= mem1702;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in10 <= mem0203;
    4'h1: pe01_in10 <= mem0303;
    4'h2: pe01_in10 <= mem0403;
    4'h3: pe01_in10 <= mem0503;
    4'h4: pe01_in10 <= mem0603;
    4'h5: pe01_in10 <= mem0703;
    4'h6: pe01_in10 <= mem0803;
    4'h7: pe01_in10 <= mem0903;
    4'h8: pe01_in10 <= mem1003;
    4'h9: pe01_in10 <= mem1103;
    4'ha: pe01_in10 <= mem1203;
    4'hb: pe01_in10 <= mem1303;
    4'hc: pe01_in10 <= mem1403;
    4'hd: pe01_in10 <= mem1503;
    4'he: pe01_in10 <= mem1603;
    4'hf: pe01_in10 <= mem1703;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in11 <= mem0204;
    4'h1: pe01_in11 <= mem0304;
    4'h2: pe01_in11 <= mem0404;
    4'h3: pe01_in11 <= mem0504;
    4'h4: pe01_in11 <= mem0604;
    4'h5: pe01_in11 <= mem0704;
    4'h6: pe01_in11 <= mem0804;
    4'h7: pe01_in11 <= mem0904;
    4'h8: pe01_in11 <= mem1004;
    4'h9: pe01_in11 <= mem1104;
    4'ha: pe01_in11 <= mem1204;
    4'hb: pe01_in11 <= mem1304;
    4'hc: pe01_in11 <= mem1404;
    4'hd: pe01_in11 <= mem1504;
    4'he: pe01_in11 <= mem1604;
    4'hf: pe01_in11 <= mem1704;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in12 <= mem0301;
    4'h1: pe01_in12 <= mem0401;
    4'h2: pe01_in12 <= mem0501;
    4'h3: pe01_in12 <= mem0601;
    4'h4: pe01_in12 <= mem0701;
    4'h5: pe01_in12 <= mem0801;
    4'h6: pe01_in12 <= mem0901;
    4'h7: pe01_in12 <= mem1001;
    4'h8: pe01_in12 <= mem1101;
    4'h9: pe01_in12 <= mem1201;
    4'ha: pe01_in12 <= mem1301;
    4'hb: pe01_in12 <= mem1401;
    4'hc: pe01_in12 <= mem1501;
    4'hd: pe01_in12 <= mem1601;
    4'he: pe01_in12 <= mem1701;
    4'hf: pe01_in12 <= mem1801;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in13 <= mem0302;
    4'h1: pe01_in13 <= mem0402;
    4'h2: pe01_in13 <= mem0502;
    4'h3: pe01_in13 <= mem0602;
    4'h4: pe01_in13 <= mem0702;
    4'h5: pe01_in13 <= mem0802;
    4'h6: pe01_in13 <= mem0902;
    4'h7: pe01_in13 <= mem1002;
    4'h8: pe01_in13 <= mem1102;
    4'h9: pe01_in13 <= mem1202;
    4'ha: pe01_in13 <= mem1302;
    4'hb: pe01_in13 <= mem1402;
    4'hc: pe01_in13 <= mem1502;
    4'hd: pe01_in13 <= mem1602;
    4'he: pe01_in13 <= mem1702;
    4'hf: pe01_in13 <= mem1802;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in14 <= mem0303;
    4'h1: pe01_in14 <= mem0403;
    4'h2: pe01_in14 <= mem0503;
    4'h3: pe01_in14 <= mem0603;
    4'h4: pe01_in14 <= mem0703;
    4'h5: pe01_in14 <= mem0803;
    4'h6: pe01_in14 <= mem0903;
    4'h7: pe01_in14 <= mem1003;
    4'h8: pe01_in14 <= mem1103;
    4'h9: pe01_in14 <= mem1203;
    4'ha: pe01_in14 <= mem1303;
    4'hb: pe01_in14 <= mem1403;
    4'hc: pe01_in14 <= mem1503;
    4'hd: pe01_in14 <= mem1603;
    4'he: pe01_in14 <= mem1703;
    4'hf: pe01_in14 <= mem1803;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe01_in15 <= mem0304;
    4'h1: pe01_in15 <= mem0404;
    4'h2: pe01_in15 <= mem0504;
    4'h3: pe01_in15 <= mem0604;
    4'h4: pe01_in15 <= mem0704;
    4'h5: pe01_in15 <= mem0804;
    4'h6: pe01_in15 <= mem0904;
    4'h7: pe01_in15 <= mem1004;
    4'h8: pe01_in15 <= mem1104;
    4'h9: pe01_in15 <= mem1204;
    4'ha: pe01_in15 <= mem1304;
    4'hb: pe01_in15 <= mem1404;
    4'hc: pe01_in15 <= mem1504;
    4'hd: pe01_in15 <= mem1604;
    4'he: pe01_in15 <= mem1704;
    4'hf: pe01_in15 <= mem1804;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in00 <= mem0002;
    4'h1: pe02_in00 <= mem0102;
    4'h2: pe02_in00 <= mem0202;
    4'h3: pe02_in00 <= mem0302;
    4'h4: pe02_in00 <= mem0402;
    4'h5: pe02_in00 <= mem0502;
    4'h6: pe02_in00 <= mem0602;
    4'h7: pe02_in00 <= mem0702;
    4'h8: pe02_in00 <= mem0802;
    4'h9: pe02_in00 <= mem0902;
    4'ha: pe02_in00 <= mem1002;
    4'hb: pe02_in00 <= mem1102;
    4'hc: pe02_in00 <= mem1202;
    4'hd: pe02_in00 <= mem1302;
    4'he: pe02_in00 <= mem1402;
    4'hf: pe02_in00 <= mem1502;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in01 <= mem0003;
    4'h1: pe02_in01 <= mem0103;
    4'h2: pe02_in01 <= mem0203;
    4'h3: pe02_in01 <= mem0303;
    4'h4: pe02_in01 <= mem0403;
    4'h5: pe02_in01 <= mem0503;
    4'h6: pe02_in01 <= mem0603;
    4'h7: pe02_in01 <= mem0703;
    4'h8: pe02_in01 <= mem0803;
    4'h9: pe02_in01 <= mem0903;
    4'ha: pe02_in01 <= mem1003;
    4'hb: pe02_in01 <= mem1103;
    4'hc: pe02_in01 <= mem1203;
    4'hd: pe02_in01 <= mem1303;
    4'he: pe02_in01 <= mem1403;
    4'hf: pe02_in01 <= mem1503;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in02 <= mem0004;
    4'h1: pe02_in02 <= mem0104;
    4'h2: pe02_in02 <= mem0204;
    4'h3: pe02_in02 <= mem0304;
    4'h4: pe02_in02 <= mem0404;
    4'h5: pe02_in02 <= mem0504;
    4'h6: pe02_in02 <= mem0604;
    4'h7: pe02_in02 <= mem0704;
    4'h8: pe02_in02 <= mem0804;
    4'h9: pe02_in02 <= mem0904;
    4'ha: pe02_in02 <= mem1004;
    4'hb: pe02_in02 <= mem1104;
    4'hc: pe02_in02 <= mem1204;
    4'hd: pe02_in02 <= mem1304;
    4'he: pe02_in02 <= mem1404;
    4'hf: pe02_in02 <= mem1504;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in03 <= mem0005;
    4'h1: pe02_in03 <= mem0105;
    4'h2: pe02_in03 <= mem0205;
    4'h3: pe02_in03 <= mem0305;
    4'h4: pe02_in03 <= mem0405;
    4'h5: pe02_in03 <= mem0505;
    4'h6: pe02_in03 <= mem0605;
    4'h7: pe02_in03 <= mem0705;
    4'h8: pe02_in03 <= mem0805;
    4'h9: pe02_in03 <= mem0905;
    4'ha: pe02_in03 <= mem1005;
    4'hb: pe02_in03 <= mem1105;
    4'hc: pe02_in03 <= mem1205;
    4'hd: pe02_in03 <= mem1305;
    4'he: pe02_in03 <= mem1405;
    4'hf: pe02_in03 <= mem1505;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in04 <= mem0102;
    4'h1: pe02_in04 <= mem0202;
    4'h2: pe02_in04 <= mem0302;
    4'h3: pe02_in04 <= mem0402;
    4'h4: pe02_in04 <= mem0502;
    4'h5: pe02_in04 <= mem0602;
    4'h6: pe02_in04 <= mem0702;
    4'h7: pe02_in04 <= mem0802;
    4'h8: pe02_in04 <= mem0902;
    4'h9: pe02_in04 <= mem1002;
    4'ha: pe02_in04 <= mem1102;
    4'hb: pe02_in04 <= mem1202;
    4'hc: pe02_in04 <= mem1302;
    4'hd: pe02_in04 <= mem1402;
    4'he: pe02_in04 <= mem1502;
    4'hf: pe02_in04 <= mem1602;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in05 <= mem0103;
    4'h1: pe02_in05 <= mem0203;
    4'h2: pe02_in05 <= mem0303;
    4'h3: pe02_in05 <= mem0403;
    4'h4: pe02_in05 <= mem0503;
    4'h5: pe02_in05 <= mem0603;
    4'h6: pe02_in05 <= mem0703;
    4'h7: pe02_in05 <= mem0803;
    4'h8: pe02_in05 <= mem0903;
    4'h9: pe02_in05 <= mem1003;
    4'ha: pe02_in05 <= mem1103;
    4'hb: pe02_in05 <= mem1203;
    4'hc: pe02_in05 <= mem1303;
    4'hd: pe02_in05 <= mem1403;
    4'he: pe02_in05 <= mem1503;
    4'hf: pe02_in05 <= mem1603;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in06 <= mem0104;
    4'h1: pe02_in06 <= mem0204;
    4'h2: pe02_in06 <= mem0304;
    4'h3: pe02_in06 <= mem0404;
    4'h4: pe02_in06 <= mem0504;
    4'h5: pe02_in06 <= mem0604;
    4'h6: pe02_in06 <= mem0704;
    4'h7: pe02_in06 <= mem0804;
    4'h8: pe02_in06 <= mem0904;
    4'h9: pe02_in06 <= mem1004;
    4'ha: pe02_in06 <= mem1104;
    4'hb: pe02_in06 <= mem1204;
    4'hc: pe02_in06 <= mem1304;
    4'hd: pe02_in06 <= mem1404;
    4'he: pe02_in06 <= mem1504;
    4'hf: pe02_in06 <= mem1604;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in07 <= mem0105;
    4'h1: pe02_in07 <= mem0205;
    4'h2: pe02_in07 <= mem0305;
    4'h3: pe02_in07 <= mem0405;
    4'h4: pe02_in07 <= mem0505;
    4'h5: pe02_in07 <= mem0605;
    4'h6: pe02_in07 <= mem0705;
    4'h7: pe02_in07 <= mem0805;
    4'h8: pe02_in07 <= mem0905;
    4'h9: pe02_in07 <= mem1005;
    4'ha: pe02_in07 <= mem1105;
    4'hb: pe02_in07 <= mem1205;
    4'hc: pe02_in07 <= mem1305;
    4'hd: pe02_in07 <= mem1405;
    4'he: pe02_in07 <= mem1505;
    4'hf: pe02_in07 <= mem1605;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in08 <= mem0202;
    4'h1: pe02_in08 <= mem0302;
    4'h2: pe02_in08 <= mem0402;
    4'h3: pe02_in08 <= mem0502;
    4'h4: pe02_in08 <= mem0602;
    4'h5: pe02_in08 <= mem0702;
    4'h6: pe02_in08 <= mem0802;
    4'h7: pe02_in08 <= mem0902;
    4'h8: pe02_in08 <= mem1002;
    4'h9: pe02_in08 <= mem1102;
    4'ha: pe02_in08 <= mem1202;
    4'hb: pe02_in08 <= mem1302;
    4'hc: pe02_in08 <= mem1402;
    4'hd: pe02_in08 <= mem1502;
    4'he: pe02_in08 <= mem1602;
    4'hf: pe02_in08 <= mem1702;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in09 <= mem0203;
    4'h1: pe02_in09 <= mem0303;
    4'h2: pe02_in09 <= mem0403;
    4'h3: pe02_in09 <= mem0503;
    4'h4: pe02_in09 <= mem0603;
    4'h5: pe02_in09 <= mem0703;
    4'h6: pe02_in09 <= mem0803;
    4'h7: pe02_in09 <= mem0903;
    4'h8: pe02_in09 <= mem1003;
    4'h9: pe02_in09 <= mem1103;
    4'ha: pe02_in09 <= mem1203;
    4'hb: pe02_in09 <= mem1303;
    4'hc: pe02_in09 <= mem1403;
    4'hd: pe02_in09 <= mem1503;
    4'he: pe02_in09 <= mem1603;
    4'hf: pe02_in09 <= mem1703;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in10 <= mem0204;
    4'h1: pe02_in10 <= mem0304;
    4'h2: pe02_in10 <= mem0404;
    4'h3: pe02_in10 <= mem0504;
    4'h4: pe02_in10 <= mem0604;
    4'h5: pe02_in10 <= mem0704;
    4'h6: pe02_in10 <= mem0804;
    4'h7: pe02_in10 <= mem0904;
    4'h8: pe02_in10 <= mem1004;
    4'h9: pe02_in10 <= mem1104;
    4'ha: pe02_in10 <= mem1204;
    4'hb: pe02_in10 <= mem1304;
    4'hc: pe02_in10 <= mem1404;
    4'hd: pe02_in10 <= mem1504;
    4'he: pe02_in10 <= mem1604;
    4'hf: pe02_in10 <= mem1704;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in11 <= mem0205;
    4'h1: pe02_in11 <= mem0305;
    4'h2: pe02_in11 <= mem0405;
    4'h3: pe02_in11 <= mem0505;
    4'h4: pe02_in11 <= mem0605;
    4'h5: pe02_in11 <= mem0705;
    4'h6: pe02_in11 <= mem0805;
    4'h7: pe02_in11 <= mem0905;
    4'h8: pe02_in11 <= mem1005;
    4'h9: pe02_in11 <= mem1105;
    4'ha: pe02_in11 <= mem1205;
    4'hb: pe02_in11 <= mem1305;
    4'hc: pe02_in11 <= mem1405;
    4'hd: pe02_in11 <= mem1505;
    4'he: pe02_in11 <= mem1605;
    4'hf: pe02_in11 <= mem1705;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in12 <= mem0302;
    4'h1: pe02_in12 <= mem0402;
    4'h2: pe02_in12 <= mem0502;
    4'h3: pe02_in12 <= mem0602;
    4'h4: pe02_in12 <= mem0702;
    4'h5: pe02_in12 <= mem0802;
    4'h6: pe02_in12 <= mem0902;
    4'h7: pe02_in12 <= mem1002;
    4'h8: pe02_in12 <= mem1102;
    4'h9: pe02_in12 <= mem1202;
    4'ha: pe02_in12 <= mem1302;
    4'hb: pe02_in12 <= mem1402;
    4'hc: pe02_in12 <= mem1502;
    4'hd: pe02_in12 <= mem1602;
    4'he: pe02_in12 <= mem1702;
    4'hf: pe02_in12 <= mem1802;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in13 <= mem0303;
    4'h1: pe02_in13 <= mem0403;
    4'h2: pe02_in13 <= mem0503;
    4'h3: pe02_in13 <= mem0603;
    4'h4: pe02_in13 <= mem0703;
    4'h5: pe02_in13 <= mem0803;
    4'h6: pe02_in13 <= mem0903;
    4'h7: pe02_in13 <= mem1003;
    4'h8: pe02_in13 <= mem1103;
    4'h9: pe02_in13 <= mem1203;
    4'ha: pe02_in13 <= mem1303;
    4'hb: pe02_in13 <= mem1403;
    4'hc: pe02_in13 <= mem1503;
    4'hd: pe02_in13 <= mem1603;
    4'he: pe02_in13 <= mem1703;
    4'hf: pe02_in13 <= mem1803;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in14 <= mem0304;
    4'h1: pe02_in14 <= mem0404;
    4'h2: pe02_in14 <= mem0504;
    4'h3: pe02_in14 <= mem0604;
    4'h4: pe02_in14 <= mem0704;
    4'h5: pe02_in14 <= mem0804;
    4'h6: pe02_in14 <= mem0904;
    4'h7: pe02_in14 <= mem1004;
    4'h8: pe02_in14 <= mem1104;
    4'h9: pe02_in14 <= mem1204;
    4'ha: pe02_in14 <= mem1304;
    4'hb: pe02_in14 <= mem1404;
    4'hc: pe02_in14 <= mem1504;
    4'hd: pe02_in14 <= mem1604;
    4'he: pe02_in14 <= mem1704;
    4'hf: pe02_in14 <= mem1804;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe02_in15 <= mem0305;
    4'h1: pe02_in15 <= mem0405;
    4'h2: pe02_in15 <= mem0505;
    4'h3: pe02_in15 <= mem0605;
    4'h4: pe02_in15 <= mem0705;
    4'h5: pe02_in15 <= mem0805;
    4'h6: pe02_in15 <= mem0905;
    4'h7: pe02_in15 <= mem1005;
    4'h8: pe02_in15 <= mem1105;
    4'h9: pe02_in15 <= mem1205;
    4'ha: pe02_in15 <= mem1305;
    4'hb: pe02_in15 <= mem1405;
    4'hc: pe02_in15 <= mem1505;
    4'hd: pe02_in15 <= mem1605;
    4'he: pe02_in15 <= mem1705;
    4'hf: pe02_in15 <= mem1805;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in00 <= mem0003;
    4'h1: pe03_in00 <= mem0103;
    4'h2: pe03_in00 <= mem0203;
    4'h3: pe03_in00 <= mem0303;
    4'h4: pe03_in00 <= mem0403;
    4'h5: pe03_in00 <= mem0503;
    4'h6: pe03_in00 <= mem0603;
    4'h7: pe03_in00 <= mem0703;
    4'h8: pe03_in00 <= mem0803;
    4'h9: pe03_in00 <= mem0903;
    4'ha: pe03_in00 <= mem1003;
    4'hb: pe03_in00 <= mem1103;
    4'hc: pe03_in00 <= mem1203;
    4'hd: pe03_in00 <= mem1303;
    4'he: pe03_in00 <= mem1403;
    4'hf: pe03_in00 <= mem1503;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in01 <= mem0004;
    4'h1: pe03_in01 <= mem0104;
    4'h2: pe03_in01 <= mem0204;
    4'h3: pe03_in01 <= mem0304;
    4'h4: pe03_in01 <= mem0404;
    4'h5: pe03_in01 <= mem0504;
    4'h6: pe03_in01 <= mem0604;
    4'h7: pe03_in01 <= mem0704;
    4'h8: pe03_in01 <= mem0804;
    4'h9: pe03_in01 <= mem0904;
    4'ha: pe03_in01 <= mem1004;
    4'hb: pe03_in01 <= mem1104;
    4'hc: pe03_in01 <= mem1204;
    4'hd: pe03_in01 <= mem1304;
    4'he: pe03_in01 <= mem1404;
    4'hf: pe03_in01 <= mem1504;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in02 <= mem0005;
    4'h1: pe03_in02 <= mem0105;
    4'h2: pe03_in02 <= mem0205;
    4'h3: pe03_in02 <= mem0305;
    4'h4: pe03_in02 <= mem0405;
    4'h5: pe03_in02 <= mem0505;
    4'h6: pe03_in02 <= mem0605;
    4'h7: pe03_in02 <= mem0705;
    4'h8: pe03_in02 <= mem0805;
    4'h9: pe03_in02 <= mem0905;
    4'ha: pe03_in02 <= mem1005;
    4'hb: pe03_in02 <= mem1105;
    4'hc: pe03_in02 <= mem1205;
    4'hd: pe03_in02 <= mem1305;
    4'he: pe03_in02 <= mem1405;
    4'hf: pe03_in02 <= mem1505;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in03 <= mem0006;
    4'h1: pe03_in03 <= mem0106;
    4'h2: pe03_in03 <= mem0206;
    4'h3: pe03_in03 <= mem0306;
    4'h4: pe03_in03 <= mem0406;
    4'h5: pe03_in03 <= mem0506;
    4'h6: pe03_in03 <= mem0606;
    4'h7: pe03_in03 <= mem0706;
    4'h8: pe03_in03 <= mem0806;
    4'h9: pe03_in03 <= mem0906;
    4'ha: pe03_in03 <= mem1006;
    4'hb: pe03_in03 <= mem1106;
    4'hc: pe03_in03 <= mem1206;
    4'hd: pe03_in03 <= mem1306;
    4'he: pe03_in03 <= mem1406;
    4'hf: pe03_in03 <= mem1506;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in04 <= mem0103;
    4'h1: pe03_in04 <= mem0203;
    4'h2: pe03_in04 <= mem0303;
    4'h3: pe03_in04 <= mem0403;
    4'h4: pe03_in04 <= mem0503;
    4'h5: pe03_in04 <= mem0603;
    4'h6: pe03_in04 <= mem0703;
    4'h7: pe03_in04 <= mem0803;
    4'h8: pe03_in04 <= mem0903;
    4'h9: pe03_in04 <= mem1003;
    4'ha: pe03_in04 <= mem1103;
    4'hb: pe03_in04 <= mem1203;
    4'hc: pe03_in04 <= mem1303;
    4'hd: pe03_in04 <= mem1403;
    4'he: pe03_in04 <= mem1503;
    4'hf: pe03_in04 <= mem1603;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in05 <= mem0104;
    4'h1: pe03_in05 <= mem0204;
    4'h2: pe03_in05 <= mem0304;
    4'h3: pe03_in05 <= mem0404;
    4'h4: pe03_in05 <= mem0504;
    4'h5: pe03_in05 <= mem0604;
    4'h6: pe03_in05 <= mem0704;
    4'h7: pe03_in05 <= mem0804;
    4'h8: pe03_in05 <= mem0904;
    4'h9: pe03_in05 <= mem1004;
    4'ha: pe03_in05 <= mem1104;
    4'hb: pe03_in05 <= mem1204;
    4'hc: pe03_in05 <= mem1304;
    4'hd: pe03_in05 <= mem1404;
    4'he: pe03_in05 <= mem1504;
    4'hf: pe03_in05 <= mem1604;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in06 <= mem0105;
    4'h1: pe03_in06 <= mem0205;
    4'h2: pe03_in06 <= mem0305;
    4'h3: pe03_in06 <= mem0405;
    4'h4: pe03_in06 <= mem0505;
    4'h5: pe03_in06 <= mem0605;
    4'h6: pe03_in06 <= mem0705;
    4'h7: pe03_in06 <= mem0805;
    4'h8: pe03_in06 <= mem0905;
    4'h9: pe03_in06 <= mem1005;
    4'ha: pe03_in06 <= mem1105;
    4'hb: pe03_in06 <= mem1205;
    4'hc: pe03_in06 <= mem1305;
    4'hd: pe03_in06 <= mem1405;
    4'he: pe03_in06 <= mem1505;
    4'hf: pe03_in06 <= mem1605;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in07 <= mem0106;
    4'h1: pe03_in07 <= mem0206;
    4'h2: pe03_in07 <= mem0306;
    4'h3: pe03_in07 <= mem0406;
    4'h4: pe03_in07 <= mem0506;
    4'h5: pe03_in07 <= mem0606;
    4'h6: pe03_in07 <= mem0706;
    4'h7: pe03_in07 <= mem0806;
    4'h8: pe03_in07 <= mem0906;
    4'h9: pe03_in07 <= mem1006;
    4'ha: pe03_in07 <= mem1106;
    4'hb: pe03_in07 <= mem1206;
    4'hc: pe03_in07 <= mem1306;
    4'hd: pe03_in07 <= mem1406;
    4'he: pe03_in07 <= mem1506;
    4'hf: pe03_in07 <= mem1606;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in08 <= mem0203;
    4'h1: pe03_in08 <= mem0303;
    4'h2: pe03_in08 <= mem0403;
    4'h3: pe03_in08 <= mem0503;
    4'h4: pe03_in08 <= mem0603;
    4'h5: pe03_in08 <= mem0703;
    4'h6: pe03_in08 <= mem0803;
    4'h7: pe03_in08 <= mem0903;
    4'h8: pe03_in08 <= mem1003;
    4'h9: pe03_in08 <= mem1103;
    4'ha: pe03_in08 <= mem1203;
    4'hb: pe03_in08 <= mem1303;
    4'hc: pe03_in08 <= mem1403;
    4'hd: pe03_in08 <= mem1503;
    4'he: pe03_in08 <= mem1603;
    4'hf: pe03_in08 <= mem1703;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in09 <= mem0204;
    4'h1: pe03_in09 <= mem0304;
    4'h2: pe03_in09 <= mem0404;
    4'h3: pe03_in09 <= mem0504;
    4'h4: pe03_in09 <= mem0604;
    4'h5: pe03_in09 <= mem0704;
    4'h6: pe03_in09 <= mem0804;
    4'h7: pe03_in09 <= mem0904;
    4'h8: pe03_in09 <= mem1004;
    4'h9: pe03_in09 <= mem1104;
    4'ha: pe03_in09 <= mem1204;
    4'hb: pe03_in09 <= mem1304;
    4'hc: pe03_in09 <= mem1404;
    4'hd: pe03_in09 <= mem1504;
    4'he: pe03_in09 <= mem1604;
    4'hf: pe03_in09 <= mem1704;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in10 <= mem0205;
    4'h1: pe03_in10 <= mem0305;
    4'h2: pe03_in10 <= mem0405;
    4'h3: pe03_in10 <= mem0505;
    4'h4: pe03_in10 <= mem0605;
    4'h5: pe03_in10 <= mem0705;
    4'h6: pe03_in10 <= mem0805;
    4'h7: pe03_in10 <= mem0905;
    4'h8: pe03_in10 <= mem1005;
    4'h9: pe03_in10 <= mem1105;
    4'ha: pe03_in10 <= mem1205;
    4'hb: pe03_in10 <= mem1305;
    4'hc: pe03_in10 <= mem1405;
    4'hd: pe03_in10 <= mem1505;
    4'he: pe03_in10 <= mem1605;
    4'hf: pe03_in10 <= mem1705;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in11 <= mem0206;
    4'h1: pe03_in11 <= mem0306;
    4'h2: pe03_in11 <= mem0406;
    4'h3: pe03_in11 <= mem0506;
    4'h4: pe03_in11 <= mem0606;
    4'h5: pe03_in11 <= mem0706;
    4'h6: pe03_in11 <= mem0806;
    4'h7: pe03_in11 <= mem0906;
    4'h8: pe03_in11 <= mem1006;
    4'h9: pe03_in11 <= mem1106;
    4'ha: pe03_in11 <= mem1206;
    4'hb: pe03_in11 <= mem1306;
    4'hc: pe03_in11 <= mem1406;
    4'hd: pe03_in11 <= mem1506;
    4'he: pe03_in11 <= mem1606;
    4'hf: pe03_in11 <= mem1706;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in12 <= mem0303;
    4'h1: pe03_in12 <= mem0403;
    4'h2: pe03_in12 <= mem0503;
    4'h3: pe03_in12 <= mem0603;
    4'h4: pe03_in12 <= mem0703;
    4'h5: pe03_in12 <= mem0803;
    4'h6: pe03_in12 <= mem0903;
    4'h7: pe03_in12 <= mem1003;
    4'h8: pe03_in12 <= mem1103;
    4'h9: pe03_in12 <= mem1203;
    4'ha: pe03_in12 <= mem1303;
    4'hb: pe03_in12 <= mem1403;
    4'hc: pe03_in12 <= mem1503;
    4'hd: pe03_in12 <= mem1603;
    4'he: pe03_in12 <= mem1703;
    4'hf: pe03_in12 <= mem1803;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in13 <= mem0304;
    4'h1: pe03_in13 <= mem0404;
    4'h2: pe03_in13 <= mem0504;
    4'h3: pe03_in13 <= mem0604;
    4'h4: pe03_in13 <= mem0704;
    4'h5: pe03_in13 <= mem0804;
    4'h6: pe03_in13 <= mem0904;
    4'h7: pe03_in13 <= mem1004;
    4'h8: pe03_in13 <= mem1104;
    4'h9: pe03_in13 <= mem1204;
    4'ha: pe03_in13 <= mem1304;
    4'hb: pe03_in13 <= mem1404;
    4'hc: pe03_in13 <= mem1504;
    4'hd: pe03_in13 <= mem1604;
    4'he: pe03_in13 <= mem1704;
    4'hf: pe03_in13 <= mem1804;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in14 <= mem0305;
    4'h1: pe03_in14 <= mem0405;
    4'h2: pe03_in14 <= mem0505;
    4'h3: pe03_in14 <= mem0605;
    4'h4: pe03_in14 <= mem0705;
    4'h5: pe03_in14 <= mem0805;
    4'h6: pe03_in14 <= mem0905;
    4'h7: pe03_in14 <= mem1005;
    4'h8: pe03_in14 <= mem1105;
    4'h9: pe03_in14 <= mem1205;
    4'ha: pe03_in14 <= mem1305;
    4'hb: pe03_in14 <= mem1405;
    4'hc: pe03_in14 <= mem1505;
    4'hd: pe03_in14 <= mem1605;
    4'he: pe03_in14 <= mem1705;
    4'hf: pe03_in14 <= mem1805;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe03_in15 <= mem0306;
    4'h1: pe03_in15 <= mem0406;
    4'h2: pe03_in15 <= mem0506;
    4'h3: pe03_in15 <= mem0606;
    4'h4: pe03_in15 <= mem0706;
    4'h5: pe03_in15 <= mem0806;
    4'h6: pe03_in15 <= mem0906;
    4'h7: pe03_in15 <= mem1006;
    4'h8: pe03_in15 <= mem1106;
    4'h9: pe03_in15 <= mem1206;
    4'ha: pe03_in15 <= mem1306;
    4'hb: pe03_in15 <= mem1406;
    4'hc: pe03_in15 <= mem1506;
    4'hd: pe03_in15 <= mem1606;
    4'he: pe03_in15 <= mem1706;
    4'hf: pe03_in15 <= mem1806;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in00 <= mem0004;
    4'h1: pe04_in00 <= mem0104;
    4'h2: pe04_in00 <= mem0204;
    4'h3: pe04_in00 <= mem0304;
    4'h4: pe04_in00 <= mem0404;
    4'h5: pe04_in00 <= mem0504;
    4'h6: pe04_in00 <= mem0604;
    4'h7: pe04_in00 <= mem0704;
    4'h8: pe04_in00 <= mem0804;
    4'h9: pe04_in00 <= mem0904;
    4'ha: pe04_in00 <= mem1004;
    4'hb: pe04_in00 <= mem1104;
    4'hc: pe04_in00 <= mem1204;
    4'hd: pe04_in00 <= mem1304;
    4'he: pe04_in00 <= mem1404;
    4'hf: pe04_in00 <= mem1504;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in01 <= mem0005;
    4'h1: pe04_in01 <= mem0105;
    4'h2: pe04_in01 <= mem0205;
    4'h3: pe04_in01 <= mem0305;
    4'h4: pe04_in01 <= mem0405;
    4'h5: pe04_in01 <= mem0505;
    4'h6: pe04_in01 <= mem0605;
    4'h7: pe04_in01 <= mem0705;
    4'h8: pe04_in01 <= mem0805;
    4'h9: pe04_in01 <= mem0905;
    4'ha: pe04_in01 <= mem1005;
    4'hb: pe04_in01 <= mem1105;
    4'hc: pe04_in01 <= mem1205;
    4'hd: pe04_in01 <= mem1305;
    4'he: pe04_in01 <= mem1405;
    4'hf: pe04_in01 <= mem1505;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in02 <= mem0006;
    4'h1: pe04_in02 <= mem0106;
    4'h2: pe04_in02 <= mem0206;
    4'h3: pe04_in02 <= mem0306;
    4'h4: pe04_in02 <= mem0406;
    4'h5: pe04_in02 <= mem0506;
    4'h6: pe04_in02 <= mem0606;
    4'h7: pe04_in02 <= mem0706;
    4'h8: pe04_in02 <= mem0806;
    4'h9: pe04_in02 <= mem0906;
    4'ha: pe04_in02 <= mem1006;
    4'hb: pe04_in02 <= mem1106;
    4'hc: pe04_in02 <= mem1206;
    4'hd: pe04_in02 <= mem1306;
    4'he: pe04_in02 <= mem1406;
    4'hf: pe04_in02 <= mem1506;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in03 <= mem0007;
    4'h1: pe04_in03 <= mem0107;
    4'h2: pe04_in03 <= mem0207;
    4'h3: pe04_in03 <= mem0307;
    4'h4: pe04_in03 <= mem0407;
    4'h5: pe04_in03 <= mem0507;
    4'h6: pe04_in03 <= mem0607;
    4'h7: pe04_in03 <= mem0707;
    4'h8: pe04_in03 <= mem0807;
    4'h9: pe04_in03 <= mem0907;
    4'ha: pe04_in03 <= mem1007;
    4'hb: pe04_in03 <= mem1107;
    4'hc: pe04_in03 <= mem1207;
    4'hd: pe04_in03 <= mem1307;
    4'he: pe04_in03 <= mem1407;
    4'hf: pe04_in03 <= mem1507;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in04 <= mem0104;
    4'h1: pe04_in04 <= mem0204;
    4'h2: pe04_in04 <= mem0304;
    4'h3: pe04_in04 <= mem0404;
    4'h4: pe04_in04 <= mem0504;
    4'h5: pe04_in04 <= mem0604;
    4'h6: pe04_in04 <= mem0704;
    4'h7: pe04_in04 <= mem0804;
    4'h8: pe04_in04 <= mem0904;
    4'h9: pe04_in04 <= mem1004;
    4'ha: pe04_in04 <= mem1104;
    4'hb: pe04_in04 <= mem1204;
    4'hc: pe04_in04 <= mem1304;
    4'hd: pe04_in04 <= mem1404;
    4'he: pe04_in04 <= mem1504;
    4'hf: pe04_in04 <= mem1604;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in05 <= mem0105;
    4'h1: pe04_in05 <= mem0205;
    4'h2: pe04_in05 <= mem0305;
    4'h3: pe04_in05 <= mem0405;
    4'h4: pe04_in05 <= mem0505;
    4'h5: pe04_in05 <= mem0605;
    4'h6: pe04_in05 <= mem0705;
    4'h7: pe04_in05 <= mem0805;
    4'h8: pe04_in05 <= mem0905;
    4'h9: pe04_in05 <= mem1005;
    4'ha: pe04_in05 <= mem1105;
    4'hb: pe04_in05 <= mem1205;
    4'hc: pe04_in05 <= mem1305;
    4'hd: pe04_in05 <= mem1405;
    4'he: pe04_in05 <= mem1505;
    4'hf: pe04_in05 <= mem1605;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in06 <= mem0106;
    4'h1: pe04_in06 <= mem0206;
    4'h2: pe04_in06 <= mem0306;
    4'h3: pe04_in06 <= mem0406;
    4'h4: pe04_in06 <= mem0506;
    4'h5: pe04_in06 <= mem0606;
    4'h6: pe04_in06 <= mem0706;
    4'h7: pe04_in06 <= mem0806;
    4'h8: pe04_in06 <= mem0906;
    4'h9: pe04_in06 <= mem1006;
    4'ha: pe04_in06 <= mem1106;
    4'hb: pe04_in06 <= mem1206;
    4'hc: pe04_in06 <= mem1306;
    4'hd: pe04_in06 <= mem1406;
    4'he: pe04_in06 <= mem1506;
    4'hf: pe04_in06 <= mem1606;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in07 <= mem0107;
    4'h1: pe04_in07 <= mem0207;
    4'h2: pe04_in07 <= mem0307;
    4'h3: pe04_in07 <= mem0407;
    4'h4: pe04_in07 <= mem0507;
    4'h5: pe04_in07 <= mem0607;
    4'h6: pe04_in07 <= mem0707;
    4'h7: pe04_in07 <= mem0807;
    4'h8: pe04_in07 <= mem0907;
    4'h9: pe04_in07 <= mem1007;
    4'ha: pe04_in07 <= mem1107;
    4'hb: pe04_in07 <= mem1207;
    4'hc: pe04_in07 <= mem1307;
    4'hd: pe04_in07 <= mem1407;
    4'he: pe04_in07 <= mem1507;
    4'hf: pe04_in07 <= mem1607;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in08 <= mem0204;
    4'h1: pe04_in08 <= mem0304;
    4'h2: pe04_in08 <= mem0404;
    4'h3: pe04_in08 <= mem0504;
    4'h4: pe04_in08 <= mem0604;
    4'h5: pe04_in08 <= mem0704;
    4'h6: pe04_in08 <= mem0804;
    4'h7: pe04_in08 <= mem0904;
    4'h8: pe04_in08 <= mem1004;
    4'h9: pe04_in08 <= mem1104;
    4'ha: pe04_in08 <= mem1204;
    4'hb: pe04_in08 <= mem1304;
    4'hc: pe04_in08 <= mem1404;
    4'hd: pe04_in08 <= mem1504;
    4'he: pe04_in08 <= mem1604;
    4'hf: pe04_in08 <= mem1704;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in09 <= mem0205;
    4'h1: pe04_in09 <= mem0305;
    4'h2: pe04_in09 <= mem0405;
    4'h3: pe04_in09 <= mem0505;
    4'h4: pe04_in09 <= mem0605;
    4'h5: pe04_in09 <= mem0705;
    4'h6: pe04_in09 <= mem0805;
    4'h7: pe04_in09 <= mem0905;
    4'h8: pe04_in09 <= mem1005;
    4'h9: pe04_in09 <= mem1105;
    4'ha: pe04_in09 <= mem1205;
    4'hb: pe04_in09 <= mem1305;
    4'hc: pe04_in09 <= mem1405;
    4'hd: pe04_in09 <= mem1505;
    4'he: pe04_in09 <= mem1605;
    4'hf: pe04_in09 <= mem1705;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in10 <= mem0206;
    4'h1: pe04_in10 <= mem0306;
    4'h2: pe04_in10 <= mem0406;
    4'h3: pe04_in10 <= mem0506;
    4'h4: pe04_in10 <= mem0606;
    4'h5: pe04_in10 <= mem0706;
    4'h6: pe04_in10 <= mem0806;
    4'h7: pe04_in10 <= mem0906;
    4'h8: pe04_in10 <= mem1006;
    4'h9: pe04_in10 <= mem1106;
    4'ha: pe04_in10 <= mem1206;
    4'hb: pe04_in10 <= mem1306;
    4'hc: pe04_in10 <= mem1406;
    4'hd: pe04_in10 <= mem1506;
    4'he: pe04_in10 <= mem1606;
    4'hf: pe04_in10 <= mem1706;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in11 <= mem0207;
    4'h1: pe04_in11 <= mem0307;
    4'h2: pe04_in11 <= mem0407;
    4'h3: pe04_in11 <= mem0507;
    4'h4: pe04_in11 <= mem0607;
    4'h5: pe04_in11 <= mem0707;
    4'h6: pe04_in11 <= mem0807;
    4'h7: pe04_in11 <= mem0907;
    4'h8: pe04_in11 <= mem1007;
    4'h9: pe04_in11 <= mem1107;
    4'ha: pe04_in11 <= mem1207;
    4'hb: pe04_in11 <= mem1307;
    4'hc: pe04_in11 <= mem1407;
    4'hd: pe04_in11 <= mem1507;
    4'he: pe04_in11 <= mem1607;
    4'hf: pe04_in11 <= mem1707;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in12 <= mem0304;
    4'h1: pe04_in12 <= mem0404;
    4'h2: pe04_in12 <= mem0504;
    4'h3: pe04_in12 <= mem0604;
    4'h4: pe04_in12 <= mem0704;
    4'h5: pe04_in12 <= mem0804;
    4'h6: pe04_in12 <= mem0904;
    4'h7: pe04_in12 <= mem1004;
    4'h8: pe04_in12 <= mem1104;
    4'h9: pe04_in12 <= mem1204;
    4'ha: pe04_in12 <= mem1304;
    4'hb: pe04_in12 <= mem1404;
    4'hc: pe04_in12 <= mem1504;
    4'hd: pe04_in12 <= mem1604;
    4'he: pe04_in12 <= mem1704;
    4'hf: pe04_in12 <= mem1804;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in13 <= mem0305;
    4'h1: pe04_in13 <= mem0405;
    4'h2: pe04_in13 <= mem0505;
    4'h3: pe04_in13 <= mem0605;
    4'h4: pe04_in13 <= mem0705;
    4'h5: pe04_in13 <= mem0805;
    4'h6: pe04_in13 <= mem0905;
    4'h7: pe04_in13 <= mem1005;
    4'h8: pe04_in13 <= mem1105;
    4'h9: pe04_in13 <= mem1205;
    4'ha: pe04_in13 <= mem1305;
    4'hb: pe04_in13 <= mem1405;
    4'hc: pe04_in13 <= mem1505;
    4'hd: pe04_in13 <= mem1605;
    4'he: pe04_in13 <= mem1705;
    4'hf: pe04_in13 <= mem1805;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in14 <= mem0306;
    4'h1: pe04_in14 <= mem0406;
    4'h2: pe04_in14 <= mem0506;
    4'h3: pe04_in14 <= mem0606;
    4'h4: pe04_in14 <= mem0706;
    4'h5: pe04_in14 <= mem0806;
    4'h6: pe04_in14 <= mem0906;
    4'h7: pe04_in14 <= mem1006;
    4'h8: pe04_in14 <= mem1106;
    4'h9: pe04_in14 <= mem1206;
    4'ha: pe04_in14 <= mem1306;
    4'hb: pe04_in14 <= mem1406;
    4'hc: pe04_in14 <= mem1506;
    4'hd: pe04_in14 <= mem1606;
    4'he: pe04_in14 <= mem1706;
    4'hf: pe04_in14 <= mem1806;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe04_in15 <= mem0307;
    4'h1: pe04_in15 <= mem0407;
    4'h2: pe04_in15 <= mem0507;
    4'h3: pe04_in15 <= mem0607;
    4'h4: pe04_in15 <= mem0707;
    4'h5: pe04_in15 <= mem0807;
    4'h6: pe04_in15 <= mem0907;
    4'h7: pe04_in15 <= mem1007;
    4'h8: pe04_in15 <= mem1107;
    4'h9: pe04_in15 <= mem1207;
    4'ha: pe04_in15 <= mem1307;
    4'hb: pe04_in15 <= mem1407;
    4'hc: pe04_in15 <= mem1507;
    4'hd: pe04_in15 <= mem1607;
    4'he: pe04_in15 <= mem1707;
    4'hf: pe04_in15 <= mem1807;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in00 <= mem0005;
    4'h1: pe05_in00 <= mem0105;
    4'h2: pe05_in00 <= mem0205;
    4'h3: pe05_in00 <= mem0305;
    4'h4: pe05_in00 <= mem0405;
    4'h5: pe05_in00 <= mem0505;
    4'h6: pe05_in00 <= mem0605;
    4'h7: pe05_in00 <= mem0705;
    4'h8: pe05_in00 <= mem0805;
    4'h9: pe05_in00 <= mem0905;
    4'ha: pe05_in00 <= mem1005;
    4'hb: pe05_in00 <= mem1105;
    4'hc: pe05_in00 <= mem1205;
    4'hd: pe05_in00 <= mem1305;
    4'he: pe05_in00 <= mem1405;
    4'hf: pe05_in00 <= mem1505;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in01 <= mem0006;
    4'h1: pe05_in01 <= mem0106;
    4'h2: pe05_in01 <= mem0206;
    4'h3: pe05_in01 <= mem0306;
    4'h4: pe05_in01 <= mem0406;
    4'h5: pe05_in01 <= mem0506;
    4'h6: pe05_in01 <= mem0606;
    4'h7: pe05_in01 <= mem0706;
    4'h8: pe05_in01 <= mem0806;
    4'h9: pe05_in01 <= mem0906;
    4'ha: pe05_in01 <= mem1006;
    4'hb: pe05_in01 <= mem1106;
    4'hc: pe05_in01 <= mem1206;
    4'hd: pe05_in01 <= mem1306;
    4'he: pe05_in01 <= mem1406;
    4'hf: pe05_in01 <= mem1506;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in02 <= mem0007;
    4'h1: pe05_in02 <= mem0107;
    4'h2: pe05_in02 <= mem0207;
    4'h3: pe05_in02 <= mem0307;
    4'h4: pe05_in02 <= mem0407;
    4'h5: pe05_in02 <= mem0507;
    4'h6: pe05_in02 <= mem0607;
    4'h7: pe05_in02 <= mem0707;
    4'h8: pe05_in02 <= mem0807;
    4'h9: pe05_in02 <= mem0907;
    4'ha: pe05_in02 <= mem1007;
    4'hb: pe05_in02 <= mem1107;
    4'hc: pe05_in02 <= mem1207;
    4'hd: pe05_in02 <= mem1307;
    4'he: pe05_in02 <= mem1407;
    4'hf: pe05_in02 <= mem1507;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in03 <= mem0008;
    4'h1: pe05_in03 <= mem0108;
    4'h2: pe05_in03 <= mem0208;
    4'h3: pe05_in03 <= mem0308;
    4'h4: pe05_in03 <= mem0408;
    4'h5: pe05_in03 <= mem0508;
    4'h6: pe05_in03 <= mem0608;
    4'h7: pe05_in03 <= mem0708;
    4'h8: pe05_in03 <= mem0808;
    4'h9: pe05_in03 <= mem0908;
    4'ha: pe05_in03 <= mem1008;
    4'hb: pe05_in03 <= mem1108;
    4'hc: pe05_in03 <= mem1208;
    4'hd: pe05_in03 <= mem1308;
    4'he: pe05_in03 <= mem1408;
    4'hf: pe05_in03 <= mem1508;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in04 <= mem0105;
    4'h1: pe05_in04 <= mem0205;
    4'h2: pe05_in04 <= mem0305;
    4'h3: pe05_in04 <= mem0405;
    4'h4: pe05_in04 <= mem0505;
    4'h5: pe05_in04 <= mem0605;
    4'h6: pe05_in04 <= mem0705;
    4'h7: pe05_in04 <= mem0805;
    4'h8: pe05_in04 <= mem0905;
    4'h9: pe05_in04 <= mem1005;
    4'ha: pe05_in04 <= mem1105;
    4'hb: pe05_in04 <= mem1205;
    4'hc: pe05_in04 <= mem1305;
    4'hd: pe05_in04 <= mem1405;
    4'he: pe05_in04 <= mem1505;
    4'hf: pe05_in04 <= mem1605;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in05 <= mem0106;
    4'h1: pe05_in05 <= mem0206;
    4'h2: pe05_in05 <= mem0306;
    4'h3: pe05_in05 <= mem0406;
    4'h4: pe05_in05 <= mem0506;
    4'h5: pe05_in05 <= mem0606;
    4'h6: pe05_in05 <= mem0706;
    4'h7: pe05_in05 <= mem0806;
    4'h8: pe05_in05 <= mem0906;
    4'h9: pe05_in05 <= mem1006;
    4'ha: pe05_in05 <= mem1106;
    4'hb: pe05_in05 <= mem1206;
    4'hc: pe05_in05 <= mem1306;
    4'hd: pe05_in05 <= mem1406;
    4'he: pe05_in05 <= mem1506;
    4'hf: pe05_in05 <= mem1606;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in06 <= mem0107;
    4'h1: pe05_in06 <= mem0207;
    4'h2: pe05_in06 <= mem0307;
    4'h3: pe05_in06 <= mem0407;
    4'h4: pe05_in06 <= mem0507;
    4'h5: pe05_in06 <= mem0607;
    4'h6: pe05_in06 <= mem0707;
    4'h7: pe05_in06 <= mem0807;
    4'h8: pe05_in06 <= mem0907;
    4'h9: pe05_in06 <= mem1007;
    4'ha: pe05_in06 <= mem1107;
    4'hb: pe05_in06 <= mem1207;
    4'hc: pe05_in06 <= mem1307;
    4'hd: pe05_in06 <= mem1407;
    4'he: pe05_in06 <= mem1507;
    4'hf: pe05_in06 <= mem1607;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in07 <= mem0108;
    4'h1: pe05_in07 <= mem0208;
    4'h2: pe05_in07 <= mem0308;
    4'h3: pe05_in07 <= mem0408;
    4'h4: pe05_in07 <= mem0508;
    4'h5: pe05_in07 <= mem0608;
    4'h6: pe05_in07 <= mem0708;
    4'h7: pe05_in07 <= mem0808;
    4'h8: pe05_in07 <= mem0908;
    4'h9: pe05_in07 <= mem1008;
    4'ha: pe05_in07 <= mem1108;
    4'hb: pe05_in07 <= mem1208;
    4'hc: pe05_in07 <= mem1308;
    4'hd: pe05_in07 <= mem1408;
    4'he: pe05_in07 <= mem1508;
    4'hf: pe05_in07 <= mem1608;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in08 <= mem0205;
    4'h1: pe05_in08 <= mem0305;
    4'h2: pe05_in08 <= mem0405;
    4'h3: pe05_in08 <= mem0505;
    4'h4: pe05_in08 <= mem0605;
    4'h5: pe05_in08 <= mem0705;
    4'h6: pe05_in08 <= mem0805;
    4'h7: pe05_in08 <= mem0905;
    4'h8: pe05_in08 <= mem1005;
    4'h9: pe05_in08 <= mem1105;
    4'ha: pe05_in08 <= mem1205;
    4'hb: pe05_in08 <= mem1305;
    4'hc: pe05_in08 <= mem1405;
    4'hd: pe05_in08 <= mem1505;
    4'he: pe05_in08 <= mem1605;
    4'hf: pe05_in08 <= mem1705;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in09 <= mem0206;
    4'h1: pe05_in09 <= mem0306;
    4'h2: pe05_in09 <= mem0406;
    4'h3: pe05_in09 <= mem0506;
    4'h4: pe05_in09 <= mem0606;
    4'h5: pe05_in09 <= mem0706;
    4'h6: pe05_in09 <= mem0806;
    4'h7: pe05_in09 <= mem0906;
    4'h8: pe05_in09 <= mem1006;
    4'h9: pe05_in09 <= mem1106;
    4'ha: pe05_in09 <= mem1206;
    4'hb: pe05_in09 <= mem1306;
    4'hc: pe05_in09 <= mem1406;
    4'hd: pe05_in09 <= mem1506;
    4'he: pe05_in09 <= mem1606;
    4'hf: pe05_in09 <= mem1706;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in10 <= mem0207;
    4'h1: pe05_in10 <= mem0307;
    4'h2: pe05_in10 <= mem0407;
    4'h3: pe05_in10 <= mem0507;
    4'h4: pe05_in10 <= mem0607;
    4'h5: pe05_in10 <= mem0707;
    4'h6: pe05_in10 <= mem0807;
    4'h7: pe05_in10 <= mem0907;
    4'h8: pe05_in10 <= mem1007;
    4'h9: pe05_in10 <= mem1107;
    4'ha: pe05_in10 <= mem1207;
    4'hb: pe05_in10 <= mem1307;
    4'hc: pe05_in10 <= mem1407;
    4'hd: pe05_in10 <= mem1507;
    4'he: pe05_in10 <= mem1607;
    4'hf: pe05_in10 <= mem1707;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in11 <= mem0208;
    4'h1: pe05_in11 <= mem0308;
    4'h2: pe05_in11 <= mem0408;
    4'h3: pe05_in11 <= mem0508;
    4'h4: pe05_in11 <= mem0608;
    4'h5: pe05_in11 <= mem0708;
    4'h6: pe05_in11 <= mem0808;
    4'h7: pe05_in11 <= mem0908;
    4'h8: pe05_in11 <= mem1008;
    4'h9: pe05_in11 <= mem1108;
    4'ha: pe05_in11 <= mem1208;
    4'hb: pe05_in11 <= mem1308;
    4'hc: pe05_in11 <= mem1408;
    4'hd: pe05_in11 <= mem1508;
    4'he: pe05_in11 <= mem1608;
    4'hf: pe05_in11 <= mem1708;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in12 <= mem0305;
    4'h1: pe05_in12 <= mem0405;
    4'h2: pe05_in12 <= mem0505;
    4'h3: pe05_in12 <= mem0605;
    4'h4: pe05_in12 <= mem0705;
    4'h5: pe05_in12 <= mem0805;
    4'h6: pe05_in12 <= mem0905;
    4'h7: pe05_in12 <= mem1005;
    4'h8: pe05_in12 <= mem1105;
    4'h9: pe05_in12 <= mem1205;
    4'ha: pe05_in12 <= mem1305;
    4'hb: pe05_in12 <= mem1405;
    4'hc: pe05_in12 <= mem1505;
    4'hd: pe05_in12 <= mem1605;
    4'he: pe05_in12 <= mem1705;
    4'hf: pe05_in12 <= mem1805;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in13 <= mem0306;
    4'h1: pe05_in13 <= mem0406;
    4'h2: pe05_in13 <= mem0506;
    4'h3: pe05_in13 <= mem0606;
    4'h4: pe05_in13 <= mem0706;
    4'h5: pe05_in13 <= mem0806;
    4'h6: pe05_in13 <= mem0906;
    4'h7: pe05_in13 <= mem1006;
    4'h8: pe05_in13 <= mem1106;
    4'h9: pe05_in13 <= mem1206;
    4'ha: pe05_in13 <= mem1306;
    4'hb: pe05_in13 <= mem1406;
    4'hc: pe05_in13 <= mem1506;
    4'hd: pe05_in13 <= mem1606;
    4'he: pe05_in13 <= mem1706;
    4'hf: pe05_in13 <= mem1806;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in14 <= mem0307;
    4'h1: pe05_in14 <= mem0407;
    4'h2: pe05_in14 <= mem0507;
    4'h3: pe05_in14 <= mem0607;
    4'h4: pe05_in14 <= mem0707;
    4'h5: pe05_in14 <= mem0807;
    4'h6: pe05_in14 <= mem0907;
    4'h7: pe05_in14 <= mem1007;
    4'h8: pe05_in14 <= mem1107;
    4'h9: pe05_in14 <= mem1207;
    4'ha: pe05_in14 <= mem1307;
    4'hb: pe05_in14 <= mem1407;
    4'hc: pe05_in14 <= mem1507;
    4'hd: pe05_in14 <= mem1607;
    4'he: pe05_in14 <= mem1707;
    4'hf: pe05_in14 <= mem1807;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe05_in15 <= mem0308;
    4'h1: pe05_in15 <= mem0408;
    4'h2: pe05_in15 <= mem0508;
    4'h3: pe05_in15 <= mem0608;
    4'h4: pe05_in15 <= mem0708;
    4'h5: pe05_in15 <= mem0808;
    4'h6: pe05_in15 <= mem0908;
    4'h7: pe05_in15 <= mem1008;
    4'h8: pe05_in15 <= mem1108;
    4'h9: pe05_in15 <= mem1208;
    4'ha: pe05_in15 <= mem1308;
    4'hb: pe05_in15 <= mem1408;
    4'hc: pe05_in15 <= mem1508;
    4'hd: pe05_in15 <= mem1608;
    4'he: pe05_in15 <= mem1708;
    4'hf: pe05_in15 <= mem1808;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in00 <= mem0006;
    4'h1: pe06_in00 <= mem0106;
    4'h2: pe06_in00 <= mem0206;
    4'h3: pe06_in00 <= mem0306;
    4'h4: pe06_in00 <= mem0406;
    4'h5: pe06_in00 <= mem0506;
    4'h6: pe06_in00 <= mem0606;
    4'h7: pe06_in00 <= mem0706;
    4'h8: pe06_in00 <= mem0806;
    4'h9: pe06_in00 <= mem0906;
    4'ha: pe06_in00 <= mem1006;
    4'hb: pe06_in00 <= mem1106;
    4'hc: pe06_in00 <= mem1206;
    4'hd: pe06_in00 <= mem1306;
    4'he: pe06_in00 <= mem1406;
    4'hf: pe06_in00 <= mem1506;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in01 <= mem0007;
    4'h1: pe06_in01 <= mem0107;
    4'h2: pe06_in01 <= mem0207;
    4'h3: pe06_in01 <= mem0307;
    4'h4: pe06_in01 <= mem0407;
    4'h5: pe06_in01 <= mem0507;
    4'h6: pe06_in01 <= mem0607;
    4'h7: pe06_in01 <= mem0707;
    4'h8: pe06_in01 <= mem0807;
    4'h9: pe06_in01 <= mem0907;
    4'ha: pe06_in01 <= mem1007;
    4'hb: pe06_in01 <= mem1107;
    4'hc: pe06_in01 <= mem1207;
    4'hd: pe06_in01 <= mem1307;
    4'he: pe06_in01 <= mem1407;
    4'hf: pe06_in01 <= mem1507;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in02 <= mem0008;
    4'h1: pe06_in02 <= mem0108;
    4'h2: pe06_in02 <= mem0208;
    4'h3: pe06_in02 <= mem0308;
    4'h4: pe06_in02 <= mem0408;
    4'h5: pe06_in02 <= mem0508;
    4'h6: pe06_in02 <= mem0608;
    4'h7: pe06_in02 <= mem0708;
    4'h8: pe06_in02 <= mem0808;
    4'h9: pe06_in02 <= mem0908;
    4'ha: pe06_in02 <= mem1008;
    4'hb: pe06_in02 <= mem1108;
    4'hc: pe06_in02 <= mem1208;
    4'hd: pe06_in02 <= mem1308;
    4'he: pe06_in02 <= mem1408;
    4'hf: pe06_in02 <= mem1508;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in03 <= mem0009;
    4'h1: pe06_in03 <= mem0109;
    4'h2: pe06_in03 <= mem0209;
    4'h3: pe06_in03 <= mem0309;
    4'h4: pe06_in03 <= mem0409;
    4'h5: pe06_in03 <= mem0509;
    4'h6: pe06_in03 <= mem0609;
    4'h7: pe06_in03 <= mem0709;
    4'h8: pe06_in03 <= mem0809;
    4'h9: pe06_in03 <= mem0909;
    4'ha: pe06_in03 <= mem1009;
    4'hb: pe06_in03 <= mem1109;
    4'hc: pe06_in03 <= mem1209;
    4'hd: pe06_in03 <= mem1309;
    4'he: pe06_in03 <= mem1409;
    4'hf: pe06_in03 <= mem1509;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in04 <= mem0106;
    4'h1: pe06_in04 <= mem0206;
    4'h2: pe06_in04 <= mem0306;
    4'h3: pe06_in04 <= mem0406;
    4'h4: pe06_in04 <= mem0506;
    4'h5: pe06_in04 <= mem0606;
    4'h6: pe06_in04 <= mem0706;
    4'h7: pe06_in04 <= mem0806;
    4'h8: pe06_in04 <= mem0906;
    4'h9: pe06_in04 <= mem1006;
    4'ha: pe06_in04 <= mem1106;
    4'hb: pe06_in04 <= mem1206;
    4'hc: pe06_in04 <= mem1306;
    4'hd: pe06_in04 <= mem1406;
    4'he: pe06_in04 <= mem1506;
    4'hf: pe06_in04 <= mem1606;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in05 <= mem0107;
    4'h1: pe06_in05 <= mem0207;
    4'h2: pe06_in05 <= mem0307;
    4'h3: pe06_in05 <= mem0407;
    4'h4: pe06_in05 <= mem0507;
    4'h5: pe06_in05 <= mem0607;
    4'h6: pe06_in05 <= mem0707;
    4'h7: pe06_in05 <= mem0807;
    4'h8: pe06_in05 <= mem0907;
    4'h9: pe06_in05 <= mem1007;
    4'ha: pe06_in05 <= mem1107;
    4'hb: pe06_in05 <= mem1207;
    4'hc: pe06_in05 <= mem1307;
    4'hd: pe06_in05 <= mem1407;
    4'he: pe06_in05 <= mem1507;
    4'hf: pe06_in05 <= mem1607;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in06 <= mem0108;
    4'h1: pe06_in06 <= mem0208;
    4'h2: pe06_in06 <= mem0308;
    4'h3: pe06_in06 <= mem0408;
    4'h4: pe06_in06 <= mem0508;
    4'h5: pe06_in06 <= mem0608;
    4'h6: pe06_in06 <= mem0708;
    4'h7: pe06_in06 <= mem0808;
    4'h8: pe06_in06 <= mem0908;
    4'h9: pe06_in06 <= mem1008;
    4'ha: pe06_in06 <= mem1108;
    4'hb: pe06_in06 <= mem1208;
    4'hc: pe06_in06 <= mem1308;
    4'hd: pe06_in06 <= mem1408;
    4'he: pe06_in06 <= mem1508;
    4'hf: pe06_in06 <= mem1608;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in07 <= mem0109;
    4'h1: pe06_in07 <= mem0209;
    4'h2: pe06_in07 <= mem0309;
    4'h3: pe06_in07 <= mem0409;
    4'h4: pe06_in07 <= mem0509;
    4'h5: pe06_in07 <= mem0609;
    4'h6: pe06_in07 <= mem0709;
    4'h7: pe06_in07 <= mem0809;
    4'h8: pe06_in07 <= mem0909;
    4'h9: pe06_in07 <= mem1009;
    4'ha: pe06_in07 <= mem1109;
    4'hb: pe06_in07 <= mem1209;
    4'hc: pe06_in07 <= mem1309;
    4'hd: pe06_in07 <= mem1409;
    4'he: pe06_in07 <= mem1509;
    4'hf: pe06_in07 <= mem1609;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in08 <= mem0206;
    4'h1: pe06_in08 <= mem0306;
    4'h2: pe06_in08 <= mem0406;
    4'h3: pe06_in08 <= mem0506;
    4'h4: pe06_in08 <= mem0606;
    4'h5: pe06_in08 <= mem0706;
    4'h6: pe06_in08 <= mem0806;
    4'h7: pe06_in08 <= mem0906;
    4'h8: pe06_in08 <= mem1006;
    4'h9: pe06_in08 <= mem1106;
    4'ha: pe06_in08 <= mem1206;
    4'hb: pe06_in08 <= mem1306;
    4'hc: pe06_in08 <= mem1406;
    4'hd: pe06_in08 <= mem1506;
    4'he: pe06_in08 <= mem1606;
    4'hf: pe06_in08 <= mem1706;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in09 <= mem0207;
    4'h1: pe06_in09 <= mem0307;
    4'h2: pe06_in09 <= mem0407;
    4'h3: pe06_in09 <= mem0507;
    4'h4: pe06_in09 <= mem0607;
    4'h5: pe06_in09 <= mem0707;
    4'h6: pe06_in09 <= mem0807;
    4'h7: pe06_in09 <= mem0907;
    4'h8: pe06_in09 <= mem1007;
    4'h9: pe06_in09 <= mem1107;
    4'ha: pe06_in09 <= mem1207;
    4'hb: pe06_in09 <= mem1307;
    4'hc: pe06_in09 <= mem1407;
    4'hd: pe06_in09 <= mem1507;
    4'he: pe06_in09 <= mem1607;
    4'hf: pe06_in09 <= mem1707;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in10 <= mem0208;
    4'h1: pe06_in10 <= mem0308;
    4'h2: pe06_in10 <= mem0408;
    4'h3: pe06_in10 <= mem0508;
    4'h4: pe06_in10 <= mem0608;
    4'h5: pe06_in10 <= mem0708;
    4'h6: pe06_in10 <= mem0808;
    4'h7: pe06_in10 <= mem0908;
    4'h8: pe06_in10 <= mem1008;
    4'h9: pe06_in10 <= mem1108;
    4'ha: pe06_in10 <= mem1208;
    4'hb: pe06_in10 <= mem1308;
    4'hc: pe06_in10 <= mem1408;
    4'hd: pe06_in10 <= mem1508;
    4'he: pe06_in10 <= mem1608;
    4'hf: pe06_in10 <= mem1708;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in11 <= mem0209;
    4'h1: pe06_in11 <= mem0309;
    4'h2: pe06_in11 <= mem0409;
    4'h3: pe06_in11 <= mem0509;
    4'h4: pe06_in11 <= mem0609;
    4'h5: pe06_in11 <= mem0709;
    4'h6: pe06_in11 <= mem0809;
    4'h7: pe06_in11 <= mem0909;
    4'h8: pe06_in11 <= mem1009;
    4'h9: pe06_in11 <= mem1109;
    4'ha: pe06_in11 <= mem1209;
    4'hb: pe06_in11 <= mem1309;
    4'hc: pe06_in11 <= mem1409;
    4'hd: pe06_in11 <= mem1509;
    4'he: pe06_in11 <= mem1609;
    4'hf: pe06_in11 <= mem1709;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in12 <= mem0306;
    4'h1: pe06_in12 <= mem0406;
    4'h2: pe06_in12 <= mem0506;
    4'h3: pe06_in12 <= mem0606;
    4'h4: pe06_in12 <= mem0706;
    4'h5: pe06_in12 <= mem0806;
    4'h6: pe06_in12 <= mem0906;
    4'h7: pe06_in12 <= mem1006;
    4'h8: pe06_in12 <= mem1106;
    4'h9: pe06_in12 <= mem1206;
    4'ha: pe06_in12 <= mem1306;
    4'hb: pe06_in12 <= mem1406;
    4'hc: pe06_in12 <= mem1506;
    4'hd: pe06_in12 <= mem1606;
    4'he: pe06_in12 <= mem1706;
    4'hf: pe06_in12 <= mem1806;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in13 <= mem0307;
    4'h1: pe06_in13 <= mem0407;
    4'h2: pe06_in13 <= mem0507;
    4'h3: pe06_in13 <= mem0607;
    4'h4: pe06_in13 <= mem0707;
    4'h5: pe06_in13 <= mem0807;
    4'h6: pe06_in13 <= mem0907;
    4'h7: pe06_in13 <= mem1007;
    4'h8: pe06_in13 <= mem1107;
    4'h9: pe06_in13 <= mem1207;
    4'ha: pe06_in13 <= mem1307;
    4'hb: pe06_in13 <= mem1407;
    4'hc: pe06_in13 <= mem1507;
    4'hd: pe06_in13 <= mem1607;
    4'he: pe06_in13 <= mem1707;
    4'hf: pe06_in13 <= mem1807;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in14 <= mem0308;
    4'h1: pe06_in14 <= mem0408;
    4'h2: pe06_in14 <= mem0508;
    4'h3: pe06_in14 <= mem0608;
    4'h4: pe06_in14 <= mem0708;
    4'h5: pe06_in14 <= mem0808;
    4'h6: pe06_in14 <= mem0908;
    4'h7: pe06_in14 <= mem1008;
    4'h8: pe06_in14 <= mem1108;
    4'h9: pe06_in14 <= mem1208;
    4'ha: pe06_in14 <= mem1308;
    4'hb: pe06_in14 <= mem1408;
    4'hc: pe06_in14 <= mem1508;
    4'hd: pe06_in14 <= mem1608;
    4'he: pe06_in14 <= mem1708;
    4'hf: pe06_in14 <= mem1808;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe06_in15 <= mem0309;
    4'h1: pe06_in15 <= mem0409;
    4'h2: pe06_in15 <= mem0509;
    4'h3: pe06_in15 <= mem0609;
    4'h4: pe06_in15 <= mem0709;
    4'h5: pe06_in15 <= mem0809;
    4'h6: pe06_in15 <= mem0909;
    4'h7: pe06_in15 <= mem1009;
    4'h8: pe06_in15 <= mem1109;
    4'h9: pe06_in15 <= mem1209;
    4'ha: pe06_in15 <= mem1309;
    4'hb: pe06_in15 <= mem1409;
    4'hc: pe06_in15 <= mem1509;
    4'hd: pe06_in15 <= mem1609;
    4'he: pe06_in15 <= mem1709;
    4'hf: pe06_in15 <= mem1809;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in00 <= mem0007;
    4'h1: pe07_in00 <= mem0107;
    4'h2: pe07_in00 <= mem0207;
    4'h3: pe07_in00 <= mem0307;
    4'h4: pe07_in00 <= mem0407;
    4'h5: pe07_in00 <= mem0507;
    4'h6: pe07_in00 <= mem0607;
    4'h7: pe07_in00 <= mem0707;
    4'h8: pe07_in00 <= mem0807;
    4'h9: pe07_in00 <= mem0907;
    4'ha: pe07_in00 <= mem1007;
    4'hb: pe07_in00 <= mem1107;
    4'hc: pe07_in00 <= mem1207;
    4'hd: pe07_in00 <= mem1307;
    4'he: pe07_in00 <= mem1407;
    4'hf: pe07_in00 <= mem1507;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in01 <= mem0008;
    4'h1: pe07_in01 <= mem0108;
    4'h2: pe07_in01 <= mem0208;
    4'h3: pe07_in01 <= mem0308;
    4'h4: pe07_in01 <= mem0408;
    4'h5: pe07_in01 <= mem0508;
    4'h6: pe07_in01 <= mem0608;
    4'h7: pe07_in01 <= mem0708;
    4'h8: pe07_in01 <= mem0808;
    4'h9: pe07_in01 <= mem0908;
    4'ha: pe07_in01 <= mem1008;
    4'hb: pe07_in01 <= mem1108;
    4'hc: pe07_in01 <= mem1208;
    4'hd: pe07_in01 <= mem1308;
    4'he: pe07_in01 <= mem1408;
    4'hf: pe07_in01 <= mem1508;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in02 <= mem0009;
    4'h1: pe07_in02 <= mem0109;
    4'h2: pe07_in02 <= mem0209;
    4'h3: pe07_in02 <= mem0309;
    4'h4: pe07_in02 <= mem0409;
    4'h5: pe07_in02 <= mem0509;
    4'h6: pe07_in02 <= mem0609;
    4'h7: pe07_in02 <= mem0709;
    4'h8: pe07_in02 <= mem0809;
    4'h9: pe07_in02 <= mem0909;
    4'ha: pe07_in02 <= mem1009;
    4'hb: pe07_in02 <= mem1109;
    4'hc: pe07_in02 <= mem1209;
    4'hd: pe07_in02 <= mem1309;
    4'he: pe07_in02 <= mem1409;
    4'hf: pe07_in02 <= mem1509;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in03 <= mem0010;
    4'h1: pe07_in03 <= mem0110;
    4'h2: pe07_in03 <= mem0210;
    4'h3: pe07_in03 <= mem0310;
    4'h4: pe07_in03 <= mem0410;
    4'h5: pe07_in03 <= mem0510;
    4'h6: pe07_in03 <= mem0610;
    4'h7: pe07_in03 <= mem0710;
    4'h8: pe07_in03 <= mem0810;
    4'h9: pe07_in03 <= mem0910;
    4'ha: pe07_in03 <= mem1010;
    4'hb: pe07_in03 <= mem1110;
    4'hc: pe07_in03 <= mem1210;
    4'hd: pe07_in03 <= mem1310;
    4'he: pe07_in03 <= mem1410;
    4'hf: pe07_in03 <= mem1510;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in04 <= mem0107;
    4'h1: pe07_in04 <= mem0207;
    4'h2: pe07_in04 <= mem0307;
    4'h3: pe07_in04 <= mem0407;
    4'h4: pe07_in04 <= mem0507;
    4'h5: pe07_in04 <= mem0607;
    4'h6: pe07_in04 <= mem0707;
    4'h7: pe07_in04 <= mem0807;
    4'h8: pe07_in04 <= mem0907;
    4'h9: pe07_in04 <= mem1007;
    4'ha: pe07_in04 <= mem1107;
    4'hb: pe07_in04 <= mem1207;
    4'hc: pe07_in04 <= mem1307;
    4'hd: pe07_in04 <= mem1407;
    4'he: pe07_in04 <= mem1507;
    4'hf: pe07_in04 <= mem1607;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in05 <= mem0108;
    4'h1: pe07_in05 <= mem0208;
    4'h2: pe07_in05 <= mem0308;
    4'h3: pe07_in05 <= mem0408;
    4'h4: pe07_in05 <= mem0508;
    4'h5: pe07_in05 <= mem0608;
    4'h6: pe07_in05 <= mem0708;
    4'h7: pe07_in05 <= mem0808;
    4'h8: pe07_in05 <= mem0908;
    4'h9: pe07_in05 <= mem1008;
    4'ha: pe07_in05 <= mem1108;
    4'hb: pe07_in05 <= mem1208;
    4'hc: pe07_in05 <= mem1308;
    4'hd: pe07_in05 <= mem1408;
    4'he: pe07_in05 <= mem1508;
    4'hf: pe07_in05 <= mem1608;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in06 <= mem0109;
    4'h1: pe07_in06 <= mem0209;
    4'h2: pe07_in06 <= mem0309;
    4'h3: pe07_in06 <= mem0409;
    4'h4: pe07_in06 <= mem0509;
    4'h5: pe07_in06 <= mem0609;
    4'h6: pe07_in06 <= mem0709;
    4'h7: pe07_in06 <= mem0809;
    4'h8: pe07_in06 <= mem0909;
    4'h9: pe07_in06 <= mem1009;
    4'ha: pe07_in06 <= mem1109;
    4'hb: pe07_in06 <= mem1209;
    4'hc: pe07_in06 <= mem1309;
    4'hd: pe07_in06 <= mem1409;
    4'he: pe07_in06 <= mem1509;
    4'hf: pe07_in06 <= mem1609;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in07 <= mem0110;
    4'h1: pe07_in07 <= mem0210;
    4'h2: pe07_in07 <= mem0310;
    4'h3: pe07_in07 <= mem0410;
    4'h4: pe07_in07 <= mem0510;
    4'h5: pe07_in07 <= mem0610;
    4'h6: pe07_in07 <= mem0710;
    4'h7: pe07_in07 <= mem0810;
    4'h8: pe07_in07 <= mem0910;
    4'h9: pe07_in07 <= mem1010;
    4'ha: pe07_in07 <= mem1110;
    4'hb: pe07_in07 <= mem1210;
    4'hc: pe07_in07 <= mem1310;
    4'hd: pe07_in07 <= mem1410;
    4'he: pe07_in07 <= mem1510;
    4'hf: pe07_in07 <= mem1610;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in08 <= mem0207;
    4'h1: pe07_in08 <= mem0307;
    4'h2: pe07_in08 <= mem0407;
    4'h3: pe07_in08 <= mem0507;
    4'h4: pe07_in08 <= mem0607;
    4'h5: pe07_in08 <= mem0707;
    4'h6: pe07_in08 <= mem0807;
    4'h7: pe07_in08 <= mem0907;
    4'h8: pe07_in08 <= mem1007;
    4'h9: pe07_in08 <= mem1107;
    4'ha: pe07_in08 <= mem1207;
    4'hb: pe07_in08 <= mem1307;
    4'hc: pe07_in08 <= mem1407;
    4'hd: pe07_in08 <= mem1507;
    4'he: pe07_in08 <= mem1607;
    4'hf: pe07_in08 <= mem1707;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in09 <= mem0208;
    4'h1: pe07_in09 <= mem0308;
    4'h2: pe07_in09 <= mem0408;
    4'h3: pe07_in09 <= mem0508;
    4'h4: pe07_in09 <= mem0608;
    4'h5: pe07_in09 <= mem0708;
    4'h6: pe07_in09 <= mem0808;
    4'h7: pe07_in09 <= mem0908;
    4'h8: pe07_in09 <= mem1008;
    4'h9: pe07_in09 <= mem1108;
    4'ha: pe07_in09 <= mem1208;
    4'hb: pe07_in09 <= mem1308;
    4'hc: pe07_in09 <= mem1408;
    4'hd: pe07_in09 <= mem1508;
    4'he: pe07_in09 <= mem1608;
    4'hf: pe07_in09 <= mem1708;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in10 <= mem0209;
    4'h1: pe07_in10 <= mem0309;
    4'h2: pe07_in10 <= mem0409;
    4'h3: pe07_in10 <= mem0509;
    4'h4: pe07_in10 <= mem0609;
    4'h5: pe07_in10 <= mem0709;
    4'h6: pe07_in10 <= mem0809;
    4'h7: pe07_in10 <= mem0909;
    4'h8: pe07_in10 <= mem1009;
    4'h9: pe07_in10 <= mem1109;
    4'ha: pe07_in10 <= mem1209;
    4'hb: pe07_in10 <= mem1309;
    4'hc: pe07_in10 <= mem1409;
    4'hd: pe07_in10 <= mem1509;
    4'he: pe07_in10 <= mem1609;
    4'hf: pe07_in10 <= mem1709;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in11 <= mem0210;
    4'h1: pe07_in11 <= mem0310;
    4'h2: pe07_in11 <= mem0410;
    4'h3: pe07_in11 <= mem0510;
    4'h4: pe07_in11 <= mem0610;
    4'h5: pe07_in11 <= mem0710;
    4'h6: pe07_in11 <= mem0810;
    4'h7: pe07_in11 <= mem0910;
    4'h8: pe07_in11 <= mem1010;
    4'h9: pe07_in11 <= mem1110;
    4'ha: pe07_in11 <= mem1210;
    4'hb: pe07_in11 <= mem1310;
    4'hc: pe07_in11 <= mem1410;
    4'hd: pe07_in11 <= mem1510;
    4'he: pe07_in11 <= mem1610;
    4'hf: pe07_in11 <= mem1710;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in12 <= mem0307;
    4'h1: pe07_in12 <= mem0407;
    4'h2: pe07_in12 <= mem0507;
    4'h3: pe07_in12 <= mem0607;
    4'h4: pe07_in12 <= mem0707;
    4'h5: pe07_in12 <= mem0807;
    4'h6: pe07_in12 <= mem0907;
    4'h7: pe07_in12 <= mem1007;
    4'h8: pe07_in12 <= mem1107;
    4'h9: pe07_in12 <= mem1207;
    4'ha: pe07_in12 <= mem1307;
    4'hb: pe07_in12 <= mem1407;
    4'hc: pe07_in12 <= mem1507;
    4'hd: pe07_in12 <= mem1607;
    4'he: pe07_in12 <= mem1707;
    4'hf: pe07_in12 <= mem1807;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in13 <= mem0308;
    4'h1: pe07_in13 <= mem0408;
    4'h2: pe07_in13 <= mem0508;
    4'h3: pe07_in13 <= mem0608;
    4'h4: pe07_in13 <= mem0708;
    4'h5: pe07_in13 <= mem0808;
    4'h6: pe07_in13 <= mem0908;
    4'h7: pe07_in13 <= mem1008;
    4'h8: pe07_in13 <= mem1108;
    4'h9: pe07_in13 <= mem1208;
    4'ha: pe07_in13 <= mem1308;
    4'hb: pe07_in13 <= mem1408;
    4'hc: pe07_in13 <= mem1508;
    4'hd: pe07_in13 <= mem1608;
    4'he: pe07_in13 <= mem1708;
    4'hf: pe07_in13 <= mem1808;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in14 <= mem0309;
    4'h1: pe07_in14 <= mem0409;
    4'h2: pe07_in14 <= mem0509;
    4'h3: pe07_in14 <= mem0609;
    4'h4: pe07_in14 <= mem0709;
    4'h5: pe07_in14 <= mem0809;
    4'h6: pe07_in14 <= mem0909;
    4'h7: pe07_in14 <= mem1009;
    4'h8: pe07_in14 <= mem1109;
    4'h9: pe07_in14 <= mem1209;
    4'ha: pe07_in14 <= mem1309;
    4'hb: pe07_in14 <= mem1409;
    4'hc: pe07_in14 <= mem1509;
    4'hd: pe07_in14 <= mem1609;
    4'he: pe07_in14 <= mem1709;
    4'hf: pe07_in14 <= mem1809;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe07_in15 <= mem0310;
    4'h1: pe07_in15 <= mem0410;
    4'h2: pe07_in15 <= mem0510;
    4'h3: pe07_in15 <= mem0610;
    4'h4: pe07_in15 <= mem0710;
    4'h5: pe07_in15 <= mem0810;
    4'h6: pe07_in15 <= mem0910;
    4'h7: pe07_in15 <= mem1010;
    4'h8: pe07_in15 <= mem1110;
    4'h9: pe07_in15 <= mem1210;
    4'ha: pe07_in15 <= mem1310;
    4'hb: pe07_in15 <= mem1410;
    4'hc: pe07_in15 <= mem1510;
    4'hd: pe07_in15 <= mem1610;
    4'he: pe07_in15 <= mem1710;
    4'hf: pe07_in15 <= mem1810;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in00 <= mem0008;
    4'h1: pe08_in00 <= mem0108;
    4'h2: pe08_in00 <= mem0208;
    4'h3: pe08_in00 <= mem0308;
    4'h4: pe08_in00 <= mem0408;
    4'h5: pe08_in00 <= mem0508;
    4'h6: pe08_in00 <= mem0608;
    4'h7: pe08_in00 <= mem0708;
    4'h8: pe08_in00 <= mem0808;
    4'h9: pe08_in00 <= mem0908;
    4'ha: pe08_in00 <= mem1008;
    4'hb: pe08_in00 <= mem1108;
    4'hc: pe08_in00 <= mem1208;
    4'hd: pe08_in00 <= mem1308;
    4'he: pe08_in00 <= mem1408;
    4'hf: pe08_in00 <= mem1508;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in01 <= mem0009;
    4'h1: pe08_in01 <= mem0109;
    4'h2: pe08_in01 <= mem0209;
    4'h3: pe08_in01 <= mem0309;
    4'h4: pe08_in01 <= mem0409;
    4'h5: pe08_in01 <= mem0509;
    4'h6: pe08_in01 <= mem0609;
    4'h7: pe08_in01 <= mem0709;
    4'h8: pe08_in01 <= mem0809;
    4'h9: pe08_in01 <= mem0909;
    4'ha: pe08_in01 <= mem1009;
    4'hb: pe08_in01 <= mem1109;
    4'hc: pe08_in01 <= mem1209;
    4'hd: pe08_in01 <= mem1309;
    4'he: pe08_in01 <= mem1409;
    4'hf: pe08_in01 <= mem1509;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in02 <= mem0010;
    4'h1: pe08_in02 <= mem0110;
    4'h2: pe08_in02 <= mem0210;
    4'h3: pe08_in02 <= mem0310;
    4'h4: pe08_in02 <= mem0410;
    4'h5: pe08_in02 <= mem0510;
    4'h6: pe08_in02 <= mem0610;
    4'h7: pe08_in02 <= mem0710;
    4'h8: pe08_in02 <= mem0810;
    4'h9: pe08_in02 <= mem0910;
    4'ha: pe08_in02 <= mem1010;
    4'hb: pe08_in02 <= mem1110;
    4'hc: pe08_in02 <= mem1210;
    4'hd: pe08_in02 <= mem1310;
    4'he: pe08_in02 <= mem1410;
    4'hf: pe08_in02 <= mem1510;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in03 <= mem0011;
    4'h1: pe08_in03 <= mem0111;
    4'h2: pe08_in03 <= mem0211;
    4'h3: pe08_in03 <= mem0311;
    4'h4: pe08_in03 <= mem0411;
    4'h5: pe08_in03 <= mem0511;
    4'h6: pe08_in03 <= mem0611;
    4'h7: pe08_in03 <= mem0711;
    4'h8: pe08_in03 <= mem0811;
    4'h9: pe08_in03 <= mem0911;
    4'ha: pe08_in03 <= mem1011;
    4'hb: pe08_in03 <= mem1111;
    4'hc: pe08_in03 <= mem1211;
    4'hd: pe08_in03 <= mem1311;
    4'he: pe08_in03 <= mem1411;
    4'hf: pe08_in03 <= mem1511;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in04 <= mem0108;
    4'h1: pe08_in04 <= mem0208;
    4'h2: pe08_in04 <= mem0308;
    4'h3: pe08_in04 <= mem0408;
    4'h4: pe08_in04 <= mem0508;
    4'h5: pe08_in04 <= mem0608;
    4'h6: pe08_in04 <= mem0708;
    4'h7: pe08_in04 <= mem0808;
    4'h8: pe08_in04 <= mem0908;
    4'h9: pe08_in04 <= mem1008;
    4'ha: pe08_in04 <= mem1108;
    4'hb: pe08_in04 <= mem1208;
    4'hc: pe08_in04 <= mem1308;
    4'hd: pe08_in04 <= mem1408;
    4'he: pe08_in04 <= mem1508;
    4'hf: pe08_in04 <= mem1608;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in05 <= mem0109;
    4'h1: pe08_in05 <= mem0209;
    4'h2: pe08_in05 <= mem0309;
    4'h3: pe08_in05 <= mem0409;
    4'h4: pe08_in05 <= mem0509;
    4'h5: pe08_in05 <= mem0609;
    4'h6: pe08_in05 <= mem0709;
    4'h7: pe08_in05 <= mem0809;
    4'h8: pe08_in05 <= mem0909;
    4'h9: pe08_in05 <= mem1009;
    4'ha: pe08_in05 <= mem1109;
    4'hb: pe08_in05 <= mem1209;
    4'hc: pe08_in05 <= mem1309;
    4'hd: pe08_in05 <= mem1409;
    4'he: pe08_in05 <= mem1509;
    4'hf: pe08_in05 <= mem1609;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in06 <= mem0110;
    4'h1: pe08_in06 <= mem0210;
    4'h2: pe08_in06 <= mem0310;
    4'h3: pe08_in06 <= mem0410;
    4'h4: pe08_in06 <= mem0510;
    4'h5: pe08_in06 <= mem0610;
    4'h6: pe08_in06 <= mem0710;
    4'h7: pe08_in06 <= mem0810;
    4'h8: pe08_in06 <= mem0910;
    4'h9: pe08_in06 <= mem1010;
    4'ha: pe08_in06 <= mem1110;
    4'hb: pe08_in06 <= mem1210;
    4'hc: pe08_in06 <= mem1310;
    4'hd: pe08_in06 <= mem1410;
    4'he: pe08_in06 <= mem1510;
    4'hf: pe08_in06 <= mem1610;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in07 <= mem0111;
    4'h1: pe08_in07 <= mem0211;
    4'h2: pe08_in07 <= mem0311;
    4'h3: pe08_in07 <= mem0411;
    4'h4: pe08_in07 <= mem0511;
    4'h5: pe08_in07 <= mem0611;
    4'h6: pe08_in07 <= mem0711;
    4'h7: pe08_in07 <= mem0811;
    4'h8: pe08_in07 <= mem0911;
    4'h9: pe08_in07 <= mem1011;
    4'ha: pe08_in07 <= mem1111;
    4'hb: pe08_in07 <= mem1211;
    4'hc: pe08_in07 <= mem1311;
    4'hd: pe08_in07 <= mem1411;
    4'he: pe08_in07 <= mem1511;
    4'hf: pe08_in07 <= mem1611;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in08 <= mem0208;
    4'h1: pe08_in08 <= mem0308;
    4'h2: pe08_in08 <= mem0408;
    4'h3: pe08_in08 <= mem0508;
    4'h4: pe08_in08 <= mem0608;
    4'h5: pe08_in08 <= mem0708;
    4'h6: pe08_in08 <= mem0808;
    4'h7: pe08_in08 <= mem0908;
    4'h8: pe08_in08 <= mem1008;
    4'h9: pe08_in08 <= mem1108;
    4'ha: pe08_in08 <= mem1208;
    4'hb: pe08_in08 <= mem1308;
    4'hc: pe08_in08 <= mem1408;
    4'hd: pe08_in08 <= mem1508;
    4'he: pe08_in08 <= mem1608;
    4'hf: pe08_in08 <= mem1708;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in09 <= mem0209;
    4'h1: pe08_in09 <= mem0309;
    4'h2: pe08_in09 <= mem0409;
    4'h3: pe08_in09 <= mem0509;
    4'h4: pe08_in09 <= mem0609;
    4'h5: pe08_in09 <= mem0709;
    4'h6: pe08_in09 <= mem0809;
    4'h7: pe08_in09 <= mem0909;
    4'h8: pe08_in09 <= mem1009;
    4'h9: pe08_in09 <= mem1109;
    4'ha: pe08_in09 <= mem1209;
    4'hb: pe08_in09 <= mem1309;
    4'hc: pe08_in09 <= mem1409;
    4'hd: pe08_in09 <= mem1509;
    4'he: pe08_in09 <= mem1609;
    4'hf: pe08_in09 <= mem1709;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in10 <= mem0210;
    4'h1: pe08_in10 <= mem0310;
    4'h2: pe08_in10 <= mem0410;
    4'h3: pe08_in10 <= mem0510;
    4'h4: pe08_in10 <= mem0610;
    4'h5: pe08_in10 <= mem0710;
    4'h6: pe08_in10 <= mem0810;
    4'h7: pe08_in10 <= mem0910;
    4'h8: pe08_in10 <= mem1010;
    4'h9: pe08_in10 <= mem1110;
    4'ha: pe08_in10 <= mem1210;
    4'hb: pe08_in10 <= mem1310;
    4'hc: pe08_in10 <= mem1410;
    4'hd: pe08_in10 <= mem1510;
    4'he: pe08_in10 <= mem1610;
    4'hf: pe08_in10 <= mem1710;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in11 <= mem0211;
    4'h1: pe08_in11 <= mem0311;
    4'h2: pe08_in11 <= mem0411;
    4'h3: pe08_in11 <= mem0511;
    4'h4: pe08_in11 <= mem0611;
    4'h5: pe08_in11 <= mem0711;
    4'h6: pe08_in11 <= mem0811;
    4'h7: pe08_in11 <= mem0911;
    4'h8: pe08_in11 <= mem1011;
    4'h9: pe08_in11 <= mem1111;
    4'ha: pe08_in11 <= mem1211;
    4'hb: pe08_in11 <= mem1311;
    4'hc: pe08_in11 <= mem1411;
    4'hd: pe08_in11 <= mem1511;
    4'he: pe08_in11 <= mem1611;
    4'hf: pe08_in11 <= mem1711;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in12 <= mem0308;
    4'h1: pe08_in12 <= mem0408;
    4'h2: pe08_in12 <= mem0508;
    4'h3: pe08_in12 <= mem0608;
    4'h4: pe08_in12 <= mem0708;
    4'h5: pe08_in12 <= mem0808;
    4'h6: pe08_in12 <= mem0908;
    4'h7: pe08_in12 <= mem1008;
    4'h8: pe08_in12 <= mem1108;
    4'h9: pe08_in12 <= mem1208;
    4'ha: pe08_in12 <= mem1308;
    4'hb: pe08_in12 <= mem1408;
    4'hc: pe08_in12 <= mem1508;
    4'hd: pe08_in12 <= mem1608;
    4'he: pe08_in12 <= mem1708;
    4'hf: pe08_in12 <= mem1808;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in13 <= mem0309;
    4'h1: pe08_in13 <= mem0409;
    4'h2: pe08_in13 <= mem0509;
    4'h3: pe08_in13 <= mem0609;
    4'h4: pe08_in13 <= mem0709;
    4'h5: pe08_in13 <= mem0809;
    4'h6: pe08_in13 <= mem0909;
    4'h7: pe08_in13 <= mem1009;
    4'h8: pe08_in13 <= mem1109;
    4'h9: pe08_in13 <= mem1209;
    4'ha: pe08_in13 <= mem1309;
    4'hb: pe08_in13 <= mem1409;
    4'hc: pe08_in13 <= mem1509;
    4'hd: pe08_in13 <= mem1609;
    4'he: pe08_in13 <= mem1709;
    4'hf: pe08_in13 <= mem1809;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in14 <= mem0310;
    4'h1: pe08_in14 <= mem0410;
    4'h2: pe08_in14 <= mem0510;
    4'h3: pe08_in14 <= mem0610;
    4'h4: pe08_in14 <= mem0710;
    4'h5: pe08_in14 <= mem0810;
    4'h6: pe08_in14 <= mem0910;
    4'h7: pe08_in14 <= mem1010;
    4'h8: pe08_in14 <= mem1110;
    4'h9: pe08_in14 <= mem1210;
    4'ha: pe08_in14 <= mem1310;
    4'hb: pe08_in14 <= mem1410;
    4'hc: pe08_in14 <= mem1510;
    4'hd: pe08_in14 <= mem1610;
    4'he: pe08_in14 <= mem1710;
    4'hf: pe08_in14 <= mem1810;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe08_in15 <= mem0311;
    4'h1: pe08_in15 <= mem0411;
    4'h2: pe08_in15 <= mem0511;
    4'h3: pe08_in15 <= mem0611;
    4'h4: pe08_in15 <= mem0711;
    4'h5: pe08_in15 <= mem0811;
    4'h6: pe08_in15 <= mem0911;
    4'h7: pe08_in15 <= mem1011;
    4'h8: pe08_in15 <= mem1111;
    4'h9: pe08_in15 <= mem1211;
    4'ha: pe08_in15 <= mem1311;
    4'hb: pe08_in15 <= mem1411;
    4'hc: pe08_in15 <= mem1511;
    4'hd: pe08_in15 <= mem1611;
    4'he: pe08_in15 <= mem1711;
    4'hf: pe08_in15 <= mem1811;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in00 <= mem0009;
    4'h1: pe09_in00 <= mem0109;
    4'h2: pe09_in00 <= mem0209;
    4'h3: pe09_in00 <= mem0309;
    4'h4: pe09_in00 <= mem0409;
    4'h5: pe09_in00 <= mem0509;
    4'h6: pe09_in00 <= mem0609;
    4'h7: pe09_in00 <= mem0709;
    4'h8: pe09_in00 <= mem0809;
    4'h9: pe09_in00 <= mem0909;
    4'ha: pe09_in00 <= mem1009;
    4'hb: pe09_in00 <= mem1109;
    4'hc: pe09_in00 <= mem1209;
    4'hd: pe09_in00 <= mem1309;
    4'he: pe09_in00 <= mem1409;
    4'hf: pe09_in00 <= mem1509;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in01 <= mem0010;
    4'h1: pe09_in01 <= mem0110;
    4'h2: pe09_in01 <= mem0210;
    4'h3: pe09_in01 <= mem0310;
    4'h4: pe09_in01 <= mem0410;
    4'h5: pe09_in01 <= mem0510;
    4'h6: pe09_in01 <= mem0610;
    4'h7: pe09_in01 <= mem0710;
    4'h8: pe09_in01 <= mem0810;
    4'h9: pe09_in01 <= mem0910;
    4'ha: pe09_in01 <= mem1010;
    4'hb: pe09_in01 <= mem1110;
    4'hc: pe09_in01 <= mem1210;
    4'hd: pe09_in01 <= mem1310;
    4'he: pe09_in01 <= mem1410;
    4'hf: pe09_in01 <= mem1510;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in02 <= mem0011;
    4'h1: pe09_in02 <= mem0111;
    4'h2: pe09_in02 <= mem0211;
    4'h3: pe09_in02 <= mem0311;
    4'h4: pe09_in02 <= mem0411;
    4'h5: pe09_in02 <= mem0511;
    4'h6: pe09_in02 <= mem0611;
    4'h7: pe09_in02 <= mem0711;
    4'h8: pe09_in02 <= mem0811;
    4'h9: pe09_in02 <= mem0911;
    4'ha: pe09_in02 <= mem1011;
    4'hb: pe09_in02 <= mem1111;
    4'hc: pe09_in02 <= mem1211;
    4'hd: pe09_in02 <= mem1311;
    4'he: pe09_in02 <= mem1411;
    4'hf: pe09_in02 <= mem1511;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in03 <= mem0012;
    4'h1: pe09_in03 <= mem0112;
    4'h2: pe09_in03 <= mem0212;
    4'h3: pe09_in03 <= mem0312;
    4'h4: pe09_in03 <= mem0412;
    4'h5: pe09_in03 <= mem0512;
    4'h6: pe09_in03 <= mem0612;
    4'h7: pe09_in03 <= mem0712;
    4'h8: pe09_in03 <= mem0812;
    4'h9: pe09_in03 <= mem0912;
    4'ha: pe09_in03 <= mem1012;
    4'hb: pe09_in03 <= mem1112;
    4'hc: pe09_in03 <= mem1212;
    4'hd: pe09_in03 <= mem1312;
    4'he: pe09_in03 <= mem1412;
    4'hf: pe09_in03 <= mem1512;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in04 <= mem0109;
    4'h1: pe09_in04 <= mem0209;
    4'h2: pe09_in04 <= mem0309;
    4'h3: pe09_in04 <= mem0409;
    4'h4: pe09_in04 <= mem0509;
    4'h5: pe09_in04 <= mem0609;
    4'h6: pe09_in04 <= mem0709;
    4'h7: pe09_in04 <= mem0809;
    4'h8: pe09_in04 <= mem0909;
    4'h9: pe09_in04 <= mem1009;
    4'ha: pe09_in04 <= mem1109;
    4'hb: pe09_in04 <= mem1209;
    4'hc: pe09_in04 <= mem1309;
    4'hd: pe09_in04 <= mem1409;
    4'he: pe09_in04 <= mem1509;
    4'hf: pe09_in04 <= mem1609;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in05 <= mem0110;
    4'h1: pe09_in05 <= mem0210;
    4'h2: pe09_in05 <= mem0310;
    4'h3: pe09_in05 <= mem0410;
    4'h4: pe09_in05 <= mem0510;
    4'h5: pe09_in05 <= mem0610;
    4'h6: pe09_in05 <= mem0710;
    4'h7: pe09_in05 <= mem0810;
    4'h8: pe09_in05 <= mem0910;
    4'h9: pe09_in05 <= mem1010;
    4'ha: pe09_in05 <= mem1110;
    4'hb: pe09_in05 <= mem1210;
    4'hc: pe09_in05 <= mem1310;
    4'hd: pe09_in05 <= mem1410;
    4'he: pe09_in05 <= mem1510;
    4'hf: pe09_in05 <= mem1610;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in06 <= mem0111;
    4'h1: pe09_in06 <= mem0211;
    4'h2: pe09_in06 <= mem0311;
    4'h3: pe09_in06 <= mem0411;
    4'h4: pe09_in06 <= mem0511;
    4'h5: pe09_in06 <= mem0611;
    4'h6: pe09_in06 <= mem0711;
    4'h7: pe09_in06 <= mem0811;
    4'h8: pe09_in06 <= mem0911;
    4'h9: pe09_in06 <= mem1011;
    4'ha: pe09_in06 <= mem1111;
    4'hb: pe09_in06 <= mem1211;
    4'hc: pe09_in06 <= mem1311;
    4'hd: pe09_in06 <= mem1411;
    4'he: pe09_in06 <= mem1511;
    4'hf: pe09_in06 <= mem1611;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in07 <= mem0112;
    4'h1: pe09_in07 <= mem0212;
    4'h2: pe09_in07 <= mem0312;
    4'h3: pe09_in07 <= mem0412;
    4'h4: pe09_in07 <= mem0512;
    4'h5: pe09_in07 <= mem0612;
    4'h6: pe09_in07 <= mem0712;
    4'h7: pe09_in07 <= mem0812;
    4'h8: pe09_in07 <= mem0912;
    4'h9: pe09_in07 <= mem1012;
    4'ha: pe09_in07 <= mem1112;
    4'hb: pe09_in07 <= mem1212;
    4'hc: pe09_in07 <= mem1312;
    4'hd: pe09_in07 <= mem1412;
    4'he: pe09_in07 <= mem1512;
    4'hf: pe09_in07 <= mem1612;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in08 <= mem0209;
    4'h1: pe09_in08 <= mem0309;
    4'h2: pe09_in08 <= mem0409;
    4'h3: pe09_in08 <= mem0509;
    4'h4: pe09_in08 <= mem0609;
    4'h5: pe09_in08 <= mem0709;
    4'h6: pe09_in08 <= mem0809;
    4'h7: pe09_in08 <= mem0909;
    4'h8: pe09_in08 <= mem1009;
    4'h9: pe09_in08 <= mem1109;
    4'ha: pe09_in08 <= mem1209;
    4'hb: pe09_in08 <= mem1309;
    4'hc: pe09_in08 <= mem1409;
    4'hd: pe09_in08 <= mem1509;
    4'he: pe09_in08 <= mem1609;
    4'hf: pe09_in08 <= mem1709;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in09 <= mem0210;
    4'h1: pe09_in09 <= mem0310;
    4'h2: pe09_in09 <= mem0410;
    4'h3: pe09_in09 <= mem0510;
    4'h4: pe09_in09 <= mem0610;
    4'h5: pe09_in09 <= mem0710;
    4'h6: pe09_in09 <= mem0810;
    4'h7: pe09_in09 <= mem0910;
    4'h8: pe09_in09 <= mem1010;
    4'h9: pe09_in09 <= mem1110;
    4'ha: pe09_in09 <= mem1210;
    4'hb: pe09_in09 <= mem1310;
    4'hc: pe09_in09 <= mem1410;
    4'hd: pe09_in09 <= mem1510;
    4'he: pe09_in09 <= mem1610;
    4'hf: pe09_in09 <= mem1710;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in10 <= mem0211;
    4'h1: pe09_in10 <= mem0311;
    4'h2: pe09_in10 <= mem0411;
    4'h3: pe09_in10 <= mem0511;
    4'h4: pe09_in10 <= mem0611;
    4'h5: pe09_in10 <= mem0711;
    4'h6: pe09_in10 <= mem0811;
    4'h7: pe09_in10 <= mem0911;
    4'h8: pe09_in10 <= mem1011;
    4'h9: pe09_in10 <= mem1111;
    4'ha: pe09_in10 <= mem1211;
    4'hb: pe09_in10 <= mem1311;
    4'hc: pe09_in10 <= mem1411;
    4'hd: pe09_in10 <= mem1511;
    4'he: pe09_in10 <= mem1611;
    4'hf: pe09_in10 <= mem1711;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in11 <= mem0212;
    4'h1: pe09_in11 <= mem0312;
    4'h2: pe09_in11 <= mem0412;
    4'h3: pe09_in11 <= mem0512;
    4'h4: pe09_in11 <= mem0612;
    4'h5: pe09_in11 <= mem0712;
    4'h6: pe09_in11 <= mem0812;
    4'h7: pe09_in11 <= mem0912;
    4'h8: pe09_in11 <= mem1012;
    4'h9: pe09_in11 <= mem1112;
    4'ha: pe09_in11 <= mem1212;
    4'hb: pe09_in11 <= mem1312;
    4'hc: pe09_in11 <= mem1412;
    4'hd: pe09_in11 <= mem1512;
    4'he: pe09_in11 <= mem1612;
    4'hf: pe09_in11 <= mem1712;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in12 <= mem0309;
    4'h1: pe09_in12 <= mem0409;
    4'h2: pe09_in12 <= mem0509;
    4'h3: pe09_in12 <= mem0609;
    4'h4: pe09_in12 <= mem0709;
    4'h5: pe09_in12 <= mem0809;
    4'h6: pe09_in12 <= mem0909;
    4'h7: pe09_in12 <= mem1009;
    4'h8: pe09_in12 <= mem1109;
    4'h9: pe09_in12 <= mem1209;
    4'ha: pe09_in12 <= mem1309;
    4'hb: pe09_in12 <= mem1409;
    4'hc: pe09_in12 <= mem1509;
    4'hd: pe09_in12 <= mem1609;
    4'he: pe09_in12 <= mem1709;
    4'hf: pe09_in12 <= mem1809;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in13 <= mem0310;
    4'h1: pe09_in13 <= mem0410;
    4'h2: pe09_in13 <= mem0510;
    4'h3: pe09_in13 <= mem0610;
    4'h4: pe09_in13 <= mem0710;
    4'h5: pe09_in13 <= mem0810;
    4'h6: pe09_in13 <= mem0910;
    4'h7: pe09_in13 <= mem1010;
    4'h8: pe09_in13 <= mem1110;
    4'h9: pe09_in13 <= mem1210;
    4'ha: pe09_in13 <= mem1310;
    4'hb: pe09_in13 <= mem1410;
    4'hc: pe09_in13 <= mem1510;
    4'hd: pe09_in13 <= mem1610;
    4'he: pe09_in13 <= mem1710;
    4'hf: pe09_in13 <= mem1810;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in14 <= mem0311;
    4'h1: pe09_in14 <= mem0411;
    4'h2: pe09_in14 <= mem0511;
    4'h3: pe09_in14 <= mem0611;
    4'h4: pe09_in14 <= mem0711;
    4'h5: pe09_in14 <= mem0811;
    4'h6: pe09_in14 <= mem0911;
    4'h7: pe09_in14 <= mem1011;
    4'h8: pe09_in14 <= mem1111;
    4'h9: pe09_in14 <= mem1211;
    4'ha: pe09_in14 <= mem1311;
    4'hb: pe09_in14 <= mem1411;
    4'hc: pe09_in14 <= mem1511;
    4'hd: pe09_in14 <= mem1611;
    4'he: pe09_in14 <= mem1711;
    4'hf: pe09_in14 <= mem1811;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe09_in15 <= mem0312;
    4'h1: pe09_in15 <= mem0412;
    4'h2: pe09_in15 <= mem0512;
    4'h3: pe09_in15 <= mem0612;
    4'h4: pe09_in15 <= mem0712;
    4'h5: pe09_in15 <= mem0812;
    4'h6: pe09_in15 <= mem0912;
    4'h7: pe09_in15 <= mem1012;
    4'h8: pe09_in15 <= mem1112;
    4'h9: pe09_in15 <= mem1212;
    4'ha: pe09_in15 <= mem1312;
    4'hb: pe09_in15 <= mem1412;
    4'hc: pe09_in15 <= mem1512;
    4'hd: pe09_in15 <= mem1612;
    4'he: pe09_in15 <= mem1712;
    4'hf: pe09_in15 <= mem1812;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in00 <= mem0010;
    4'h1: pe10_in00 <= mem0110;
    4'h2: pe10_in00 <= mem0210;
    4'h3: pe10_in00 <= mem0310;
    4'h4: pe10_in00 <= mem0410;
    4'h5: pe10_in00 <= mem0510;
    4'h6: pe10_in00 <= mem0610;
    4'h7: pe10_in00 <= mem0710;
    4'h8: pe10_in00 <= mem0810;
    4'h9: pe10_in00 <= mem0910;
    4'ha: pe10_in00 <= mem1010;
    4'hb: pe10_in00 <= mem1110;
    4'hc: pe10_in00 <= mem1210;
    4'hd: pe10_in00 <= mem1310;
    4'he: pe10_in00 <= mem1410;
    4'hf: pe10_in00 <= mem1510;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in01 <= mem0011;
    4'h1: pe10_in01 <= mem0111;
    4'h2: pe10_in01 <= mem0211;
    4'h3: pe10_in01 <= mem0311;
    4'h4: pe10_in01 <= mem0411;
    4'h5: pe10_in01 <= mem0511;
    4'h6: pe10_in01 <= mem0611;
    4'h7: pe10_in01 <= mem0711;
    4'h8: pe10_in01 <= mem0811;
    4'h9: pe10_in01 <= mem0911;
    4'ha: pe10_in01 <= mem1011;
    4'hb: pe10_in01 <= mem1111;
    4'hc: pe10_in01 <= mem1211;
    4'hd: pe10_in01 <= mem1311;
    4'he: pe10_in01 <= mem1411;
    4'hf: pe10_in01 <= mem1511;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in02 <= mem0012;
    4'h1: pe10_in02 <= mem0112;
    4'h2: pe10_in02 <= mem0212;
    4'h3: pe10_in02 <= mem0312;
    4'h4: pe10_in02 <= mem0412;
    4'h5: pe10_in02 <= mem0512;
    4'h6: pe10_in02 <= mem0612;
    4'h7: pe10_in02 <= mem0712;
    4'h8: pe10_in02 <= mem0812;
    4'h9: pe10_in02 <= mem0912;
    4'ha: pe10_in02 <= mem1012;
    4'hb: pe10_in02 <= mem1112;
    4'hc: pe10_in02 <= mem1212;
    4'hd: pe10_in02 <= mem1312;
    4'he: pe10_in02 <= mem1412;
    4'hf: pe10_in02 <= mem1512;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in03 <= mem0013;
    4'h1: pe10_in03 <= mem0113;
    4'h2: pe10_in03 <= mem0213;
    4'h3: pe10_in03 <= mem0313;
    4'h4: pe10_in03 <= mem0413;
    4'h5: pe10_in03 <= mem0513;
    4'h6: pe10_in03 <= mem0613;
    4'h7: pe10_in03 <= mem0713;
    4'h8: pe10_in03 <= mem0813;
    4'h9: pe10_in03 <= mem0913;
    4'ha: pe10_in03 <= mem1013;
    4'hb: pe10_in03 <= mem1113;
    4'hc: pe10_in03 <= mem1213;
    4'hd: pe10_in03 <= mem1313;
    4'he: pe10_in03 <= mem1413;
    4'hf: pe10_in03 <= mem1513;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in04 <= mem0110;
    4'h1: pe10_in04 <= mem0210;
    4'h2: pe10_in04 <= mem0310;
    4'h3: pe10_in04 <= mem0410;
    4'h4: pe10_in04 <= mem0510;
    4'h5: pe10_in04 <= mem0610;
    4'h6: pe10_in04 <= mem0710;
    4'h7: pe10_in04 <= mem0810;
    4'h8: pe10_in04 <= mem0910;
    4'h9: pe10_in04 <= mem1010;
    4'ha: pe10_in04 <= mem1110;
    4'hb: pe10_in04 <= mem1210;
    4'hc: pe10_in04 <= mem1310;
    4'hd: pe10_in04 <= mem1410;
    4'he: pe10_in04 <= mem1510;
    4'hf: pe10_in04 <= mem1610;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in05 <= mem0111;
    4'h1: pe10_in05 <= mem0211;
    4'h2: pe10_in05 <= mem0311;
    4'h3: pe10_in05 <= mem0411;
    4'h4: pe10_in05 <= mem0511;
    4'h5: pe10_in05 <= mem0611;
    4'h6: pe10_in05 <= mem0711;
    4'h7: pe10_in05 <= mem0811;
    4'h8: pe10_in05 <= mem0911;
    4'h9: pe10_in05 <= mem1011;
    4'ha: pe10_in05 <= mem1111;
    4'hb: pe10_in05 <= mem1211;
    4'hc: pe10_in05 <= mem1311;
    4'hd: pe10_in05 <= mem1411;
    4'he: pe10_in05 <= mem1511;
    4'hf: pe10_in05 <= mem1611;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in06 <= mem0112;
    4'h1: pe10_in06 <= mem0212;
    4'h2: pe10_in06 <= mem0312;
    4'h3: pe10_in06 <= mem0412;
    4'h4: pe10_in06 <= mem0512;
    4'h5: pe10_in06 <= mem0612;
    4'h6: pe10_in06 <= mem0712;
    4'h7: pe10_in06 <= mem0812;
    4'h8: pe10_in06 <= mem0912;
    4'h9: pe10_in06 <= mem1012;
    4'ha: pe10_in06 <= mem1112;
    4'hb: pe10_in06 <= mem1212;
    4'hc: pe10_in06 <= mem1312;
    4'hd: pe10_in06 <= mem1412;
    4'he: pe10_in06 <= mem1512;
    4'hf: pe10_in06 <= mem1612;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in07 <= mem0113;
    4'h1: pe10_in07 <= mem0213;
    4'h2: pe10_in07 <= mem0313;
    4'h3: pe10_in07 <= mem0413;
    4'h4: pe10_in07 <= mem0513;
    4'h5: pe10_in07 <= mem0613;
    4'h6: pe10_in07 <= mem0713;
    4'h7: pe10_in07 <= mem0813;
    4'h8: pe10_in07 <= mem0913;
    4'h9: pe10_in07 <= mem1013;
    4'ha: pe10_in07 <= mem1113;
    4'hb: pe10_in07 <= mem1213;
    4'hc: pe10_in07 <= mem1313;
    4'hd: pe10_in07 <= mem1413;
    4'he: pe10_in07 <= mem1513;
    4'hf: pe10_in07 <= mem1613;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in08 <= mem0210;
    4'h1: pe10_in08 <= mem0310;
    4'h2: pe10_in08 <= mem0410;
    4'h3: pe10_in08 <= mem0510;
    4'h4: pe10_in08 <= mem0610;
    4'h5: pe10_in08 <= mem0710;
    4'h6: pe10_in08 <= mem0810;
    4'h7: pe10_in08 <= mem0910;
    4'h8: pe10_in08 <= mem1010;
    4'h9: pe10_in08 <= mem1110;
    4'ha: pe10_in08 <= mem1210;
    4'hb: pe10_in08 <= mem1310;
    4'hc: pe10_in08 <= mem1410;
    4'hd: pe10_in08 <= mem1510;
    4'he: pe10_in08 <= mem1610;
    4'hf: pe10_in08 <= mem1710;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in09 <= mem0211;
    4'h1: pe10_in09 <= mem0311;
    4'h2: pe10_in09 <= mem0411;
    4'h3: pe10_in09 <= mem0511;
    4'h4: pe10_in09 <= mem0611;
    4'h5: pe10_in09 <= mem0711;
    4'h6: pe10_in09 <= mem0811;
    4'h7: pe10_in09 <= mem0911;
    4'h8: pe10_in09 <= mem1011;
    4'h9: pe10_in09 <= mem1111;
    4'ha: pe10_in09 <= mem1211;
    4'hb: pe10_in09 <= mem1311;
    4'hc: pe10_in09 <= mem1411;
    4'hd: pe10_in09 <= mem1511;
    4'he: pe10_in09 <= mem1611;
    4'hf: pe10_in09 <= mem1711;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in10 <= mem0212;
    4'h1: pe10_in10 <= mem0312;
    4'h2: pe10_in10 <= mem0412;
    4'h3: pe10_in10 <= mem0512;
    4'h4: pe10_in10 <= mem0612;
    4'h5: pe10_in10 <= mem0712;
    4'h6: pe10_in10 <= mem0812;
    4'h7: pe10_in10 <= mem0912;
    4'h8: pe10_in10 <= mem1012;
    4'h9: pe10_in10 <= mem1112;
    4'ha: pe10_in10 <= mem1212;
    4'hb: pe10_in10 <= mem1312;
    4'hc: pe10_in10 <= mem1412;
    4'hd: pe10_in10 <= mem1512;
    4'he: pe10_in10 <= mem1612;
    4'hf: pe10_in10 <= mem1712;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in11 <= mem0213;
    4'h1: pe10_in11 <= mem0313;
    4'h2: pe10_in11 <= mem0413;
    4'h3: pe10_in11 <= mem0513;
    4'h4: pe10_in11 <= mem0613;
    4'h5: pe10_in11 <= mem0713;
    4'h6: pe10_in11 <= mem0813;
    4'h7: pe10_in11 <= mem0913;
    4'h8: pe10_in11 <= mem1013;
    4'h9: pe10_in11 <= mem1113;
    4'ha: pe10_in11 <= mem1213;
    4'hb: pe10_in11 <= mem1313;
    4'hc: pe10_in11 <= mem1413;
    4'hd: pe10_in11 <= mem1513;
    4'he: pe10_in11 <= mem1613;
    4'hf: pe10_in11 <= mem1713;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in12 <= mem0310;
    4'h1: pe10_in12 <= mem0410;
    4'h2: pe10_in12 <= mem0510;
    4'h3: pe10_in12 <= mem0610;
    4'h4: pe10_in12 <= mem0710;
    4'h5: pe10_in12 <= mem0810;
    4'h6: pe10_in12 <= mem0910;
    4'h7: pe10_in12 <= mem1010;
    4'h8: pe10_in12 <= mem1110;
    4'h9: pe10_in12 <= mem1210;
    4'ha: pe10_in12 <= mem1310;
    4'hb: pe10_in12 <= mem1410;
    4'hc: pe10_in12 <= mem1510;
    4'hd: pe10_in12 <= mem1610;
    4'he: pe10_in12 <= mem1710;
    4'hf: pe10_in12 <= mem1810;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in13 <= mem0311;
    4'h1: pe10_in13 <= mem0411;
    4'h2: pe10_in13 <= mem0511;
    4'h3: pe10_in13 <= mem0611;
    4'h4: pe10_in13 <= mem0711;
    4'h5: pe10_in13 <= mem0811;
    4'h6: pe10_in13 <= mem0911;
    4'h7: pe10_in13 <= mem1011;
    4'h8: pe10_in13 <= mem1111;
    4'h9: pe10_in13 <= mem1211;
    4'ha: pe10_in13 <= mem1311;
    4'hb: pe10_in13 <= mem1411;
    4'hc: pe10_in13 <= mem1511;
    4'hd: pe10_in13 <= mem1611;
    4'he: pe10_in13 <= mem1711;
    4'hf: pe10_in13 <= mem1811;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in14 <= mem0312;
    4'h1: pe10_in14 <= mem0412;
    4'h2: pe10_in14 <= mem0512;
    4'h3: pe10_in14 <= mem0612;
    4'h4: pe10_in14 <= mem0712;
    4'h5: pe10_in14 <= mem0812;
    4'h6: pe10_in14 <= mem0912;
    4'h7: pe10_in14 <= mem1012;
    4'h8: pe10_in14 <= mem1112;
    4'h9: pe10_in14 <= mem1212;
    4'ha: pe10_in14 <= mem1312;
    4'hb: pe10_in14 <= mem1412;
    4'hc: pe10_in14 <= mem1512;
    4'hd: pe10_in14 <= mem1612;
    4'he: pe10_in14 <= mem1712;
    4'hf: pe10_in14 <= mem1812;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe10_in15 <= mem0313;
    4'h1: pe10_in15 <= mem0413;
    4'h2: pe10_in15 <= mem0513;
    4'h3: pe10_in15 <= mem0613;
    4'h4: pe10_in15 <= mem0713;
    4'h5: pe10_in15 <= mem0813;
    4'h6: pe10_in15 <= mem0913;
    4'h7: pe10_in15 <= mem1013;
    4'h8: pe10_in15 <= mem1113;
    4'h9: pe10_in15 <= mem1213;
    4'ha: pe10_in15 <= mem1313;
    4'hb: pe10_in15 <= mem1413;
    4'hc: pe10_in15 <= mem1513;
    4'hd: pe10_in15 <= mem1613;
    4'he: pe10_in15 <= mem1713;
    4'hf: pe10_in15 <= mem1813;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in00 <= mem0011;
    4'h1: pe11_in00 <= mem0111;
    4'h2: pe11_in00 <= mem0211;
    4'h3: pe11_in00 <= mem0311;
    4'h4: pe11_in00 <= mem0411;
    4'h5: pe11_in00 <= mem0511;
    4'h6: pe11_in00 <= mem0611;
    4'h7: pe11_in00 <= mem0711;
    4'h8: pe11_in00 <= mem0811;
    4'h9: pe11_in00 <= mem0911;
    4'ha: pe11_in00 <= mem1011;
    4'hb: pe11_in00 <= mem1111;
    4'hc: pe11_in00 <= mem1211;
    4'hd: pe11_in00 <= mem1311;
    4'he: pe11_in00 <= mem1411;
    4'hf: pe11_in00 <= mem1511;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in01 <= mem0012;
    4'h1: pe11_in01 <= mem0112;
    4'h2: pe11_in01 <= mem0212;
    4'h3: pe11_in01 <= mem0312;
    4'h4: pe11_in01 <= mem0412;
    4'h5: pe11_in01 <= mem0512;
    4'h6: pe11_in01 <= mem0612;
    4'h7: pe11_in01 <= mem0712;
    4'h8: pe11_in01 <= mem0812;
    4'h9: pe11_in01 <= mem0912;
    4'ha: pe11_in01 <= mem1012;
    4'hb: pe11_in01 <= mem1112;
    4'hc: pe11_in01 <= mem1212;
    4'hd: pe11_in01 <= mem1312;
    4'he: pe11_in01 <= mem1412;
    4'hf: pe11_in01 <= mem1512;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in02 <= mem0013;
    4'h1: pe11_in02 <= mem0113;
    4'h2: pe11_in02 <= mem0213;
    4'h3: pe11_in02 <= mem0313;
    4'h4: pe11_in02 <= mem0413;
    4'h5: pe11_in02 <= mem0513;
    4'h6: pe11_in02 <= mem0613;
    4'h7: pe11_in02 <= mem0713;
    4'h8: pe11_in02 <= mem0813;
    4'h9: pe11_in02 <= mem0913;
    4'ha: pe11_in02 <= mem1013;
    4'hb: pe11_in02 <= mem1113;
    4'hc: pe11_in02 <= mem1213;
    4'hd: pe11_in02 <= mem1313;
    4'he: pe11_in02 <= mem1413;
    4'hf: pe11_in02 <= mem1513;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in03 <= mem0014;
    4'h1: pe11_in03 <= mem0114;
    4'h2: pe11_in03 <= mem0214;
    4'h3: pe11_in03 <= mem0314;
    4'h4: pe11_in03 <= mem0414;
    4'h5: pe11_in03 <= mem0514;
    4'h6: pe11_in03 <= mem0614;
    4'h7: pe11_in03 <= mem0714;
    4'h8: pe11_in03 <= mem0814;
    4'h9: pe11_in03 <= mem0914;
    4'ha: pe11_in03 <= mem1014;
    4'hb: pe11_in03 <= mem1114;
    4'hc: pe11_in03 <= mem1214;
    4'hd: pe11_in03 <= mem1314;
    4'he: pe11_in03 <= mem1414;
    4'hf: pe11_in03 <= mem1514;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in04 <= mem0111;
    4'h1: pe11_in04 <= mem0211;
    4'h2: pe11_in04 <= mem0311;
    4'h3: pe11_in04 <= mem0411;
    4'h4: pe11_in04 <= mem0511;
    4'h5: pe11_in04 <= mem0611;
    4'h6: pe11_in04 <= mem0711;
    4'h7: pe11_in04 <= mem0811;
    4'h8: pe11_in04 <= mem0911;
    4'h9: pe11_in04 <= mem1011;
    4'ha: pe11_in04 <= mem1111;
    4'hb: pe11_in04 <= mem1211;
    4'hc: pe11_in04 <= mem1311;
    4'hd: pe11_in04 <= mem1411;
    4'he: pe11_in04 <= mem1511;
    4'hf: pe11_in04 <= mem1611;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in05 <= mem0112;
    4'h1: pe11_in05 <= mem0212;
    4'h2: pe11_in05 <= mem0312;
    4'h3: pe11_in05 <= mem0412;
    4'h4: pe11_in05 <= mem0512;
    4'h5: pe11_in05 <= mem0612;
    4'h6: pe11_in05 <= mem0712;
    4'h7: pe11_in05 <= mem0812;
    4'h8: pe11_in05 <= mem0912;
    4'h9: pe11_in05 <= mem1012;
    4'ha: pe11_in05 <= mem1112;
    4'hb: pe11_in05 <= mem1212;
    4'hc: pe11_in05 <= mem1312;
    4'hd: pe11_in05 <= mem1412;
    4'he: pe11_in05 <= mem1512;
    4'hf: pe11_in05 <= mem1612;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in06 <= mem0113;
    4'h1: pe11_in06 <= mem0213;
    4'h2: pe11_in06 <= mem0313;
    4'h3: pe11_in06 <= mem0413;
    4'h4: pe11_in06 <= mem0513;
    4'h5: pe11_in06 <= mem0613;
    4'h6: pe11_in06 <= mem0713;
    4'h7: pe11_in06 <= mem0813;
    4'h8: pe11_in06 <= mem0913;
    4'h9: pe11_in06 <= mem1013;
    4'ha: pe11_in06 <= mem1113;
    4'hb: pe11_in06 <= mem1213;
    4'hc: pe11_in06 <= mem1313;
    4'hd: pe11_in06 <= mem1413;
    4'he: pe11_in06 <= mem1513;
    4'hf: pe11_in06 <= mem1613;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in07 <= mem0114;
    4'h1: pe11_in07 <= mem0214;
    4'h2: pe11_in07 <= mem0314;
    4'h3: pe11_in07 <= mem0414;
    4'h4: pe11_in07 <= mem0514;
    4'h5: pe11_in07 <= mem0614;
    4'h6: pe11_in07 <= mem0714;
    4'h7: pe11_in07 <= mem0814;
    4'h8: pe11_in07 <= mem0914;
    4'h9: pe11_in07 <= mem1014;
    4'ha: pe11_in07 <= mem1114;
    4'hb: pe11_in07 <= mem1214;
    4'hc: pe11_in07 <= mem1314;
    4'hd: pe11_in07 <= mem1414;
    4'he: pe11_in07 <= mem1514;
    4'hf: pe11_in07 <= mem1614;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in08 <= mem0211;
    4'h1: pe11_in08 <= mem0311;
    4'h2: pe11_in08 <= mem0411;
    4'h3: pe11_in08 <= mem0511;
    4'h4: pe11_in08 <= mem0611;
    4'h5: pe11_in08 <= mem0711;
    4'h6: pe11_in08 <= mem0811;
    4'h7: pe11_in08 <= mem0911;
    4'h8: pe11_in08 <= mem1011;
    4'h9: pe11_in08 <= mem1111;
    4'ha: pe11_in08 <= mem1211;
    4'hb: pe11_in08 <= mem1311;
    4'hc: pe11_in08 <= mem1411;
    4'hd: pe11_in08 <= mem1511;
    4'he: pe11_in08 <= mem1611;
    4'hf: pe11_in08 <= mem1711;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in09 <= mem0212;
    4'h1: pe11_in09 <= mem0312;
    4'h2: pe11_in09 <= mem0412;
    4'h3: pe11_in09 <= mem0512;
    4'h4: pe11_in09 <= mem0612;
    4'h5: pe11_in09 <= mem0712;
    4'h6: pe11_in09 <= mem0812;
    4'h7: pe11_in09 <= mem0912;
    4'h8: pe11_in09 <= mem1012;
    4'h9: pe11_in09 <= mem1112;
    4'ha: pe11_in09 <= mem1212;
    4'hb: pe11_in09 <= mem1312;
    4'hc: pe11_in09 <= mem1412;
    4'hd: pe11_in09 <= mem1512;
    4'he: pe11_in09 <= mem1612;
    4'hf: pe11_in09 <= mem1712;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in10 <= mem0213;
    4'h1: pe11_in10 <= mem0313;
    4'h2: pe11_in10 <= mem0413;
    4'h3: pe11_in10 <= mem0513;
    4'h4: pe11_in10 <= mem0613;
    4'h5: pe11_in10 <= mem0713;
    4'h6: pe11_in10 <= mem0813;
    4'h7: pe11_in10 <= mem0913;
    4'h8: pe11_in10 <= mem1013;
    4'h9: pe11_in10 <= mem1113;
    4'ha: pe11_in10 <= mem1213;
    4'hb: pe11_in10 <= mem1313;
    4'hc: pe11_in10 <= mem1413;
    4'hd: pe11_in10 <= mem1513;
    4'he: pe11_in10 <= mem1613;
    4'hf: pe11_in10 <= mem1713;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in11 <= mem0214;
    4'h1: pe11_in11 <= mem0314;
    4'h2: pe11_in11 <= mem0414;
    4'h3: pe11_in11 <= mem0514;
    4'h4: pe11_in11 <= mem0614;
    4'h5: pe11_in11 <= mem0714;
    4'h6: pe11_in11 <= mem0814;
    4'h7: pe11_in11 <= mem0914;
    4'h8: pe11_in11 <= mem1014;
    4'h9: pe11_in11 <= mem1114;
    4'ha: pe11_in11 <= mem1214;
    4'hb: pe11_in11 <= mem1314;
    4'hc: pe11_in11 <= mem1414;
    4'hd: pe11_in11 <= mem1514;
    4'he: pe11_in11 <= mem1614;
    4'hf: pe11_in11 <= mem1714;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in12 <= mem0311;
    4'h1: pe11_in12 <= mem0411;
    4'h2: pe11_in12 <= mem0511;
    4'h3: pe11_in12 <= mem0611;
    4'h4: pe11_in12 <= mem0711;
    4'h5: pe11_in12 <= mem0811;
    4'h6: pe11_in12 <= mem0911;
    4'h7: pe11_in12 <= mem1011;
    4'h8: pe11_in12 <= mem1111;
    4'h9: pe11_in12 <= mem1211;
    4'ha: pe11_in12 <= mem1311;
    4'hb: pe11_in12 <= mem1411;
    4'hc: pe11_in12 <= mem1511;
    4'hd: pe11_in12 <= mem1611;
    4'he: pe11_in12 <= mem1711;
    4'hf: pe11_in12 <= mem1811;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in13 <= mem0312;
    4'h1: pe11_in13 <= mem0412;
    4'h2: pe11_in13 <= mem0512;
    4'h3: pe11_in13 <= mem0612;
    4'h4: pe11_in13 <= mem0712;
    4'h5: pe11_in13 <= mem0812;
    4'h6: pe11_in13 <= mem0912;
    4'h7: pe11_in13 <= mem1012;
    4'h8: pe11_in13 <= mem1112;
    4'h9: pe11_in13 <= mem1212;
    4'ha: pe11_in13 <= mem1312;
    4'hb: pe11_in13 <= mem1412;
    4'hc: pe11_in13 <= mem1512;
    4'hd: pe11_in13 <= mem1612;
    4'he: pe11_in13 <= mem1712;
    4'hf: pe11_in13 <= mem1812;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in14 <= mem0313;
    4'h1: pe11_in14 <= mem0413;
    4'h2: pe11_in14 <= mem0513;
    4'h3: pe11_in14 <= mem0613;
    4'h4: pe11_in14 <= mem0713;
    4'h5: pe11_in14 <= mem0813;
    4'h6: pe11_in14 <= mem0913;
    4'h7: pe11_in14 <= mem1013;
    4'h8: pe11_in14 <= mem1113;
    4'h9: pe11_in14 <= mem1213;
    4'ha: pe11_in14 <= mem1313;
    4'hb: pe11_in14 <= mem1413;
    4'hc: pe11_in14 <= mem1513;
    4'hd: pe11_in14 <= mem1613;
    4'he: pe11_in14 <= mem1713;
    4'hf: pe11_in14 <= mem1813;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe11_in15 <= mem0314;
    4'h1: pe11_in15 <= mem0414;
    4'h2: pe11_in15 <= mem0514;
    4'h3: pe11_in15 <= mem0614;
    4'h4: pe11_in15 <= mem0714;
    4'h5: pe11_in15 <= mem0814;
    4'h6: pe11_in15 <= mem0914;
    4'h7: pe11_in15 <= mem1014;
    4'h8: pe11_in15 <= mem1114;
    4'h9: pe11_in15 <= mem1214;
    4'ha: pe11_in15 <= mem1314;
    4'hb: pe11_in15 <= mem1414;
    4'hc: pe11_in15 <= mem1514;
    4'hd: pe11_in15 <= mem1614;
    4'he: pe11_in15 <= mem1714;
    4'hf: pe11_in15 <= mem1814;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in00 <= mem0012;
    4'h1: pe12_in00 <= mem0112;
    4'h2: pe12_in00 <= mem0212;
    4'h3: pe12_in00 <= mem0312;
    4'h4: pe12_in00 <= mem0412;
    4'h5: pe12_in00 <= mem0512;
    4'h6: pe12_in00 <= mem0612;
    4'h7: pe12_in00 <= mem0712;
    4'h8: pe12_in00 <= mem0812;
    4'h9: pe12_in00 <= mem0912;
    4'ha: pe12_in00 <= mem1012;
    4'hb: pe12_in00 <= mem1112;
    4'hc: pe12_in00 <= mem1212;
    4'hd: pe12_in00 <= mem1312;
    4'he: pe12_in00 <= mem1412;
    4'hf: pe12_in00 <= mem1512;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in01 <= mem0013;
    4'h1: pe12_in01 <= mem0113;
    4'h2: pe12_in01 <= mem0213;
    4'h3: pe12_in01 <= mem0313;
    4'h4: pe12_in01 <= mem0413;
    4'h5: pe12_in01 <= mem0513;
    4'h6: pe12_in01 <= mem0613;
    4'h7: pe12_in01 <= mem0713;
    4'h8: pe12_in01 <= mem0813;
    4'h9: pe12_in01 <= mem0913;
    4'ha: pe12_in01 <= mem1013;
    4'hb: pe12_in01 <= mem1113;
    4'hc: pe12_in01 <= mem1213;
    4'hd: pe12_in01 <= mem1313;
    4'he: pe12_in01 <= mem1413;
    4'hf: pe12_in01 <= mem1513;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in02 <= mem0014;
    4'h1: pe12_in02 <= mem0114;
    4'h2: pe12_in02 <= mem0214;
    4'h3: pe12_in02 <= mem0314;
    4'h4: pe12_in02 <= mem0414;
    4'h5: pe12_in02 <= mem0514;
    4'h6: pe12_in02 <= mem0614;
    4'h7: pe12_in02 <= mem0714;
    4'h8: pe12_in02 <= mem0814;
    4'h9: pe12_in02 <= mem0914;
    4'ha: pe12_in02 <= mem1014;
    4'hb: pe12_in02 <= mem1114;
    4'hc: pe12_in02 <= mem1214;
    4'hd: pe12_in02 <= mem1314;
    4'he: pe12_in02 <= mem1414;
    4'hf: pe12_in02 <= mem1514;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in03 <= mem0015;
    4'h1: pe12_in03 <= mem0115;
    4'h2: pe12_in03 <= mem0215;
    4'h3: pe12_in03 <= mem0315;
    4'h4: pe12_in03 <= mem0415;
    4'h5: pe12_in03 <= mem0515;
    4'h6: pe12_in03 <= mem0615;
    4'h7: pe12_in03 <= mem0715;
    4'h8: pe12_in03 <= mem0815;
    4'h9: pe12_in03 <= mem0915;
    4'ha: pe12_in03 <= mem1015;
    4'hb: pe12_in03 <= mem1115;
    4'hc: pe12_in03 <= mem1215;
    4'hd: pe12_in03 <= mem1315;
    4'he: pe12_in03 <= mem1415;
    4'hf: pe12_in03 <= mem1515;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in04 <= mem0112;
    4'h1: pe12_in04 <= mem0212;
    4'h2: pe12_in04 <= mem0312;
    4'h3: pe12_in04 <= mem0412;
    4'h4: pe12_in04 <= mem0512;
    4'h5: pe12_in04 <= mem0612;
    4'h6: pe12_in04 <= mem0712;
    4'h7: pe12_in04 <= mem0812;
    4'h8: pe12_in04 <= mem0912;
    4'h9: pe12_in04 <= mem1012;
    4'ha: pe12_in04 <= mem1112;
    4'hb: pe12_in04 <= mem1212;
    4'hc: pe12_in04 <= mem1312;
    4'hd: pe12_in04 <= mem1412;
    4'he: pe12_in04 <= mem1512;
    4'hf: pe12_in04 <= mem1612;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in05 <= mem0113;
    4'h1: pe12_in05 <= mem0213;
    4'h2: pe12_in05 <= mem0313;
    4'h3: pe12_in05 <= mem0413;
    4'h4: pe12_in05 <= mem0513;
    4'h5: pe12_in05 <= mem0613;
    4'h6: pe12_in05 <= mem0713;
    4'h7: pe12_in05 <= mem0813;
    4'h8: pe12_in05 <= mem0913;
    4'h9: pe12_in05 <= mem1013;
    4'ha: pe12_in05 <= mem1113;
    4'hb: pe12_in05 <= mem1213;
    4'hc: pe12_in05 <= mem1313;
    4'hd: pe12_in05 <= mem1413;
    4'he: pe12_in05 <= mem1513;
    4'hf: pe12_in05 <= mem1613;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in06 <= mem0114;
    4'h1: pe12_in06 <= mem0214;
    4'h2: pe12_in06 <= mem0314;
    4'h3: pe12_in06 <= mem0414;
    4'h4: pe12_in06 <= mem0514;
    4'h5: pe12_in06 <= mem0614;
    4'h6: pe12_in06 <= mem0714;
    4'h7: pe12_in06 <= mem0814;
    4'h8: pe12_in06 <= mem0914;
    4'h9: pe12_in06 <= mem1014;
    4'ha: pe12_in06 <= mem1114;
    4'hb: pe12_in06 <= mem1214;
    4'hc: pe12_in06 <= mem1314;
    4'hd: pe12_in06 <= mem1414;
    4'he: pe12_in06 <= mem1514;
    4'hf: pe12_in06 <= mem1614;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in07 <= mem0115;
    4'h1: pe12_in07 <= mem0215;
    4'h2: pe12_in07 <= mem0315;
    4'h3: pe12_in07 <= mem0415;
    4'h4: pe12_in07 <= mem0515;
    4'h5: pe12_in07 <= mem0615;
    4'h6: pe12_in07 <= mem0715;
    4'h7: pe12_in07 <= mem0815;
    4'h8: pe12_in07 <= mem0915;
    4'h9: pe12_in07 <= mem1015;
    4'ha: pe12_in07 <= mem1115;
    4'hb: pe12_in07 <= mem1215;
    4'hc: pe12_in07 <= mem1315;
    4'hd: pe12_in07 <= mem1415;
    4'he: pe12_in07 <= mem1515;
    4'hf: pe12_in07 <= mem1615;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in08 <= mem0212;
    4'h1: pe12_in08 <= mem0312;
    4'h2: pe12_in08 <= mem0412;
    4'h3: pe12_in08 <= mem0512;
    4'h4: pe12_in08 <= mem0612;
    4'h5: pe12_in08 <= mem0712;
    4'h6: pe12_in08 <= mem0812;
    4'h7: pe12_in08 <= mem0912;
    4'h8: pe12_in08 <= mem1012;
    4'h9: pe12_in08 <= mem1112;
    4'ha: pe12_in08 <= mem1212;
    4'hb: pe12_in08 <= mem1312;
    4'hc: pe12_in08 <= mem1412;
    4'hd: pe12_in08 <= mem1512;
    4'he: pe12_in08 <= mem1612;
    4'hf: pe12_in08 <= mem1712;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in09 <= mem0213;
    4'h1: pe12_in09 <= mem0313;
    4'h2: pe12_in09 <= mem0413;
    4'h3: pe12_in09 <= mem0513;
    4'h4: pe12_in09 <= mem0613;
    4'h5: pe12_in09 <= mem0713;
    4'h6: pe12_in09 <= mem0813;
    4'h7: pe12_in09 <= mem0913;
    4'h8: pe12_in09 <= mem1013;
    4'h9: pe12_in09 <= mem1113;
    4'ha: pe12_in09 <= mem1213;
    4'hb: pe12_in09 <= mem1313;
    4'hc: pe12_in09 <= mem1413;
    4'hd: pe12_in09 <= mem1513;
    4'he: pe12_in09 <= mem1613;
    4'hf: pe12_in09 <= mem1713;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in10 <= mem0214;
    4'h1: pe12_in10 <= mem0314;
    4'h2: pe12_in10 <= mem0414;
    4'h3: pe12_in10 <= mem0514;
    4'h4: pe12_in10 <= mem0614;
    4'h5: pe12_in10 <= mem0714;
    4'h6: pe12_in10 <= mem0814;
    4'h7: pe12_in10 <= mem0914;
    4'h8: pe12_in10 <= mem1014;
    4'h9: pe12_in10 <= mem1114;
    4'ha: pe12_in10 <= mem1214;
    4'hb: pe12_in10 <= mem1314;
    4'hc: pe12_in10 <= mem1414;
    4'hd: pe12_in10 <= mem1514;
    4'he: pe12_in10 <= mem1614;
    4'hf: pe12_in10 <= mem1714;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in11 <= mem0215;
    4'h1: pe12_in11 <= mem0315;
    4'h2: pe12_in11 <= mem0415;
    4'h3: pe12_in11 <= mem0515;
    4'h4: pe12_in11 <= mem0615;
    4'h5: pe12_in11 <= mem0715;
    4'h6: pe12_in11 <= mem0815;
    4'h7: pe12_in11 <= mem0915;
    4'h8: pe12_in11 <= mem1015;
    4'h9: pe12_in11 <= mem1115;
    4'ha: pe12_in11 <= mem1215;
    4'hb: pe12_in11 <= mem1315;
    4'hc: pe12_in11 <= mem1415;
    4'hd: pe12_in11 <= mem1515;
    4'he: pe12_in11 <= mem1615;
    4'hf: pe12_in11 <= mem1715;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in12 <= mem0312;
    4'h1: pe12_in12 <= mem0412;
    4'h2: pe12_in12 <= mem0512;
    4'h3: pe12_in12 <= mem0612;
    4'h4: pe12_in12 <= mem0712;
    4'h5: pe12_in12 <= mem0812;
    4'h6: pe12_in12 <= mem0912;
    4'h7: pe12_in12 <= mem1012;
    4'h8: pe12_in12 <= mem1112;
    4'h9: pe12_in12 <= mem1212;
    4'ha: pe12_in12 <= mem1312;
    4'hb: pe12_in12 <= mem1412;
    4'hc: pe12_in12 <= mem1512;
    4'hd: pe12_in12 <= mem1612;
    4'he: pe12_in12 <= mem1712;
    4'hf: pe12_in12 <= mem1812;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in13 <= mem0313;
    4'h1: pe12_in13 <= mem0413;
    4'h2: pe12_in13 <= mem0513;
    4'h3: pe12_in13 <= mem0613;
    4'h4: pe12_in13 <= mem0713;
    4'h5: pe12_in13 <= mem0813;
    4'h6: pe12_in13 <= mem0913;
    4'h7: pe12_in13 <= mem1013;
    4'h8: pe12_in13 <= mem1113;
    4'h9: pe12_in13 <= mem1213;
    4'ha: pe12_in13 <= mem1313;
    4'hb: pe12_in13 <= mem1413;
    4'hc: pe12_in13 <= mem1513;
    4'hd: pe12_in13 <= mem1613;
    4'he: pe12_in13 <= mem1713;
    4'hf: pe12_in13 <= mem1813;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in14 <= mem0314;
    4'h1: pe12_in14 <= mem0414;
    4'h2: pe12_in14 <= mem0514;
    4'h3: pe12_in14 <= mem0614;
    4'h4: pe12_in14 <= mem0714;
    4'h5: pe12_in14 <= mem0814;
    4'h6: pe12_in14 <= mem0914;
    4'h7: pe12_in14 <= mem1014;
    4'h8: pe12_in14 <= mem1114;
    4'h9: pe12_in14 <= mem1214;
    4'ha: pe12_in14 <= mem1314;
    4'hb: pe12_in14 <= mem1414;
    4'hc: pe12_in14 <= mem1514;
    4'hd: pe12_in14 <= mem1614;
    4'he: pe12_in14 <= mem1714;
    4'hf: pe12_in14 <= mem1814;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe12_in15 <= mem0315;
    4'h1: pe12_in15 <= mem0415;
    4'h2: pe12_in15 <= mem0515;
    4'h3: pe12_in15 <= mem0615;
    4'h4: pe12_in15 <= mem0715;
    4'h5: pe12_in15 <= mem0815;
    4'h6: pe12_in15 <= mem0915;
    4'h7: pe12_in15 <= mem1015;
    4'h8: pe12_in15 <= mem1115;
    4'h9: pe12_in15 <= mem1215;
    4'ha: pe12_in15 <= mem1315;
    4'hb: pe12_in15 <= mem1415;
    4'hc: pe12_in15 <= mem1515;
    4'hd: pe12_in15 <= mem1615;
    4'he: pe12_in15 <= mem1715;
    4'hf: pe12_in15 <= mem1815;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in00 <= mem0013;
    4'h1: pe13_in00 <= mem0113;
    4'h2: pe13_in00 <= mem0213;
    4'h3: pe13_in00 <= mem0313;
    4'h4: pe13_in00 <= mem0413;
    4'h5: pe13_in00 <= mem0513;
    4'h6: pe13_in00 <= mem0613;
    4'h7: pe13_in00 <= mem0713;
    4'h8: pe13_in00 <= mem0813;
    4'h9: pe13_in00 <= mem0913;
    4'ha: pe13_in00 <= mem1013;
    4'hb: pe13_in00 <= mem1113;
    4'hc: pe13_in00 <= mem1213;
    4'hd: pe13_in00 <= mem1313;
    4'he: pe13_in00 <= mem1413;
    4'hf: pe13_in00 <= mem1513;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in01 <= mem0014;
    4'h1: pe13_in01 <= mem0114;
    4'h2: pe13_in01 <= mem0214;
    4'h3: pe13_in01 <= mem0314;
    4'h4: pe13_in01 <= mem0414;
    4'h5: pe13_in01 <= mem0514;
    4'h6: pe13_in01 <= mem0614;
    4'h7: pe13_in01 <= mem0714;
    4'h8: pe13_in01 <= mem0814;
    4'h9: pe13_in01 <= mem0914;
    4'ha: pe13_in01 <= mem1014;
    4'hb: pe13_in01 <= mem1114;
    4'hc: pe13_in01 <= mem1214;
    4'hd: pe13_in01 <= mem1314;
    4'he: pe13_in01 <= mem1414;
    4'hf: pe13_in01 <= mem1514;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in02 <= mem0015;
    4'h1: pe13_in02 <= mem0115;
    4'h2: pe13_in02 <= mem0215;
    4'h3: pe13_in02 <= mem0315;
    4'h4: pe13_in02 <= mem0415;
    4'h5: pe13_in02 <= mem0515;
    4'h6: pe13_in02 <= mem0615;
    4'h7: pe13_in02 <= mem0715;
    4'h8: pe13_in02 <= mem0815;
    4'h9: pe13_in02 <= mem0915;
    4'ha: pe13_in02 <= mem1015;
    4'hb: pe13_in02 <= mem1115;
    4'hc: pe13_in02 <= mem1215;
    4'hd: pe13_in02 <= mem1315;
    4'he: pe13_in02 <= mem1415;
    4'hf: pe13_in02 <= mem1515;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in03 <= mem0016;
    4'h1: pe13_in03 <= mem0116;
    4'h2: pe13_in03 <= mem0216;
    4'h3: pe13_in03 <= mem0316;
    4'h4: pe13_in03 <= mem0416;
    4'h5: pe13_in03 <= mem0516;
    4'h6: pe13_in03 <= mem0616;
    4'h7: pe13_in03 <= mem0716;
    4'h8: pe13_in03 <= mem0816;
    4'h9: pe13_in03 <= mem0916;
    4'ha: pe13_in03 <= mem1016;
    4'hb: pe13_in03 <= mem1116;
    4'hc: pe13_in03 <= mem1216;
    4'hd: pe13_in03 <= mem1316;
    4'he: pe13_in03 <= mem1416;
    4'hf: pe13_in03 <= mem1516;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in04 <= mem0113;
    4'h1: pe13_in04 <= mem0213;
    4'h2: pe13_in04 <= mem0313;
    4'h3: pe13_in04 <= mem0413;
    4'h4: pe13_in04 <= mem0513;
    4'h5: pe13_in04 <= mem0613;
    4'h6: pe13_in04 <= mem0713;
    4'h7: pe13_in04 <= mem0813;
    4'h8: pe13_in04 <= mem0913;
    4'h9: pe13_in04 <= mem1013;
    4'ha: pe13_in04 <= mem1113;
    4'hb: pe13_in04 <= mem1213;
    4'hc: pe13_in04 <= mem1313;
    4'hd: pe13_in04 <= mem1413;
    4'he: pe13_in04 <= mem1513;
    4'hf: pe13_in04 <= mem1613;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in05 <= mem0114;
    4'h1: pe13_in05 <= mem0214;
    4'h2: pe13_in05 <= mem0314;
    4'h3: pe13_in05 <= mem0414;
    4'h4: pe13_in05 <= mem0514;
    4'h5: pe13_in05 <= mem0614;
    4'h6: pe13_in05 <= mem0714;
    4'h7: pe13_in05 <= mem0814;
    4'h8: pe13_in05 <= mem0914;
    4'h9: pe13_in05 <= mem1014;
    4'ha: pe13_in05 <= mem1114;
    4'hb: pe13_in05 <= mem1214;
    4'hc: pe13_in05 <= mem1314;
    4'hd: pe13_in05 <= mem1414;
    4'he: pe13_in05 <= mem1514;
    4'hf: pe13_in05 <= mem1614;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in06 <= mem0115;
    4'h1: pe13_in06 <= mem0215;
    4'h2: pe13_in06 <= mem0315;
    4'h3: pe13_in06 <= mem0415;
    4'h4: pe13_in06 <= mem0515;
    4'h5: pe13_in06 <= mem0615;
    4'h6: pe13_in06 <= mem0715;
    4'h7: pe13_in06 <= mem0815;
    4'h8: pe13_in06 <= mem0915;
    4'h9: pe13_in06 <= mem1015;
    4'ha: pe13_in06 <= mem1115;
    4'hb: pe13_in06 <= mem1215;
    4'hc: pe13_in06 <= mem1315;
    4'hd: pe13_in06 <= mem1415;
    4'he: pe13_in06 <= mem1515;
    4'hf: pe13_in06 <= mem1615;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in07 <= mem0116;
    4'h1: pe13_in07 <= mem0216;
    4'h2: pe13_in07 <= mem0316;
    4'h3: pe13_in07 <= mem0416;
    4'h4: pe13_in07 <= mem0516;
    4'h5: pe13_in07 <= mem0616;
    4'h6: pe13_in07 <= mem0716;
    4'h7: pe13_in07 <= mem0816;
    4'h8: pe13_in07 <= mem0916;
    4'h9: pe13_in07 <= mem1016;
    4'ha: pe13_in07 <= mem1116;
    4'hb: pe13_in07 <= mem1216;
    4'hc: pe13_in07 <= mem1316;
    4'hd: pe13_in07 <= mem1416;
    4'he: pe13_in07 <= mem1516;
    4'hf: pe13_in07 <= mem1616;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in08 <= mem0213;
    4'h1: pe13_in08 <= mem0313;
    4'h2: pe13_in08 <= mem0413;
    4'h3: pe13_in08 <= mem0513;
    4'h4: pe13_in08 <= mem0613;
    4'h5: pe13_in08 <= mem0713;
    4'h6: pe13_in08 <= mem0813;
    4'h7: pe13_in08 <= mem0913;
    4'h8: pe13_in08 <= mem1013;
    4'h9: pe13_in08 <= mem1113;
    4'ha: pe13_in08 <= mem1213;
    4'hb: pe13_in08 <= mem1313;
    4'hc: pe13_in08 <= mem1413;
    4'hd: pe13_in08 <= mem1513;
    4'he: pe13_in08 <= mem1613;
    4'hf: pe13_in08 <= mem1713;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in09 <= mem0214;
    4'h1: pe13_in09 <= mem0314;
    4'h2: pe13_in09 <= mem0414;
    4'h3: pe13_in09 <= mem0514;
    4'h4: pe13_in09 <= mem0614;
    4'h5: pe13_in09 <= mem0714;
    4'h6: pe13_in09 <= mem0814;
    4'h7: pe13_in09 <= mem0914;
    4'h8: pe13_in09 <= mem1014;
    4'h9: pe13_in09 <= mem1114;
    4'ha: pe13_in09 <= mem1214;
    4'hb: pe13_in09 <= mem1314;
    4'hc: pe13_in09 <= mem1414;
    4'hd: pe13_in09 <= mem1514;
    4'he: pe13_in09 <= mem1614;
    4'hf: pe13_in09 <= mem1714;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in10 <= mem0215;
    4'h1: pe13_in10 <= mem0315;
    4'h2: pe13_in10 <= mem0415;
    4'h3: pe13_in10 <= mem0515;
    4'h4: pe13_in10 <= mem0615;
    4'h5: pe13_in10 <= mem0715;
    4'h6: pe13_in10 <= mem0815;
    4'h7: pe13_in10 <= mem0915;
    4'h8: pe13_in10 <= mem1015;
    4'h9: pe13_in10 <= mem1115;
    4'ha: pe13_in10 <= mem1215;
    4'hb: pe13_in10 <= mem1315;
    4'hc: pe13_in10 <= mem1415;
    4'hd: pe13_in10 <= mem1515;
    4'he: pe13_in10 <= mem1615;
    4'hf: pe13_in10 <= mem1715;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in11 <= mem0216;
    4'h1: pe13_in11 <= mem0316;
    4'h2: pe13_in11 <= mem0416;
    4'h3: pe13_in11 <= mem0516;
    4'h4: pe13_in11 <= mem0616;
    4'h5: pe13_in11 <= mem0716;
    4'h6: pe13_in11 <= mem0816;
    4'h7: pe13_in11 <= mem0916;
    4'h8: pe13_in11 <= mem1016;
    4'h9: pe13_in11 <= mem1116;
    4'ha: pe13_in11 <= mem1216;
    4'hb: pe13_in11 <= mem1316;
    4'hc: pe13_in11 <= mem1416;
    4'hd: pe13_in11 <= mem1516;
    4'he: pe13_in11 <= mem1616;
    4'hf: pe13_in11 <= mem1716;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in12 <= mem0313;
    4'h1: pe13_in12 <= mem0413;
    4'h2: pe13_in12 <= mem0513;
    4'h3: pe13_in12 <= mem0613;
    4'h4: pe13_in12 <= mem0713;
    4'h5: pe13_in12 <= mem0813;
    4'h6: pe13_in12 <= mem0913;
    4'h7: pe13_in12 <= mem1013;
    4'h8: pe13_in12 <= mem1113;
    4'h9: pe13_in12 <= mem1213;
    4'ha: pe13_in12 <= mem1313;
    4'hb: pe13_in12 <= mem1413;
    4'hc: pe13_in12 <= mem1513;
    4'hd: pe13_in12 <= mem1613;
    4'he: pe13_in12 <= mem1713;
    4'hf: pe13_in12 <= mem1813;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in13 <= mem0314;
    4'h1: pe13_in13 <= mem0414;
    4'h2: pe13_in13 <= mem0514;
    4'h3: pe13_in13 <= mem0614;
    4'h4: pe13_in13 <= mem0714;
    4'h5: pe13_in13 <= mem0814;
    4'h6: pe13_in13 <= mem0914;
    4'h7: pe13_in13 <= mem1014;
    4'h8: pe13_in13 <= mem1114;
    4'h9: pe13_in13 <= mem1214;
    4'ha: pe13_in13 <= mem1314;
    4'hb: pe13_in13 <= mem1414;
    4'hc: pe13_in13 <= mem1514;
    4'hd: pe13_in13 <= mem1614;
    4'he: pe13_in13 <= mem1714;
    4'hf: pe13_in13 <= mem1814;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in14 <= mem0315;
    4'h1: pe13_in14 <= mem0415;
    4'h2: pe13_in14 <= mem0515;
    4'h3: pe13_in14 <= mem0615;
    4'h4: pe13_in14 <= mem0715;
    4'h5: pe13_in14 <= mem0815;
    4'h6: pe13_in14 <= mem0915;
    4'h7: pe13_in14 <= mem1015;
    4'h8: pe13_in14 <= mem1115;
    4'h9: pe13_in14 <= mem1215;
    4'ha: pe13_in14 <= mem1315;
    4'hb: pe13_in14 <= mem1415;
    4'hc: pe13_in14 <= mem1515;
    4'hd: pe13_in14 <= mem1615;
    4'he: pe13_in14 <= mem1715;
    4'hf: pe13_in14 <= mem1815;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe13_in15 <= mem0316;
    4'h1: pe13_in15 <= mem0416;
    4'h2: pe13_in15 <= mem0516;
    4'h3: pe13_in15 <= mem0616;
    4'h4: pe13_in15 <= mem0716;
    4'h5: pe13_in15 <= mem0816;
    4'h6: pe13_in15 <= mem0916;
    4'h7: pe13_in15 <= mem1016;
    4'h8: pe13_in15 <= mem1116;
    4'h9: pe13_in15 <= mem1216;
    4'ha: pe13_in15 <= mem1316;
    4'hb: pe13_in15 <= mem1416;
    4'hc: pe13_in15 <= mem1516;
    4'hd: pe13_in15 <= mem1616;
    4'he: pe13_in15 <= mem1716;
    4'hf: pe13_in15 <= mem1816;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in00 <= mem0014;
    4'h1: pe14_in00 <= mem0114;
    4'h2: pe14_in00 <= mem0214;
    4'h3: pe14_in00 <= mem0314;
    4'h4: pe14_in00 <= mem0414;
    4'h5: pe14_in00 <= mem0514;
    4'h6: pe14_in00 <= mem0614;
    4'h7: pe14_in00 <= mem0714;
    4'h8: pe14_in00 <= mem0814;
    4'h9: pe14_in00 <= mem0914;
    4'ha: pe14_in00 <= mem1014;
    4'hb: pe14_in00 <= mem1114;
    4'hc: pe14_in00 <= mem1214;
    4'hd: pe14_in00 <= mem1314;
    4'he: pe14_in00 <= mem1414;
    4'hf: pe14_in00 <= mem1514;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in01 <= mem0015;
    4'h1: pe14_in01 <= mem0115;
    4'h2: pe14_in01 <= mem0215;
    4'h3: pe14_in01 <= mem0315;
    4'h4: pe14_in01 <= mem0415;
    4'h5: pe14_in01 <= mem0515;
    4'h6: pe14_in01 <= mem0615;
    4'h7: pe14_in01 <= mem0715;
    4'h8: pe14_in01 <= mem0815;
    4'h9: pe14_in01 <= mem0915;
    4'ha: pe14_in01 <= mem1015;
    4'hb: pe14_in01 <= mem1115;
    4'hc: pe14_in01 <= mem1215;
    4'hd: pe14_in01 <= mem1315;
    4'he: pe14_in01 <= mem1415;
    4'hf: pe14_in01 <= mem1515;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in02 <= mem0016;
    4'h1: pe14_in02 <= mem0116;
    4'h2: pe14_in02 <= mem0216;
    4'h3: pe14_in02 <= mem0316;
    4'h4: pe14_in02 <= mem0416;
    4'h5: pe14_in02 <= mem0516;
    4'h6: pe14_in02 <= mem0616;
    4'h7: pe14_in02 <= mem0716;
    4'h8: pe14_in02 <= mem0816;
    4'h9: pe14_in02 <= mem0916;
    4'ha: pe14_in02 <= mem1016;
    4'hb: pe14_in02 <= mem1116;
    4'hc: pe14_in02 <= mem1216;
    4'hd: pe14_in02 <= mem1316;
    4'he: pe14_in02 <= mem1416;
    4'hf: pe14_in02 <= mem1516;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in03 <= mem0017;
    4'h1: pe14_in03 <= mem0117;
    4'h2: pe14_in03 <= mem0217;
    4'h3: pe14_in03 <= mem0317;
    4'h4: pe14_in03 <= mem0417;
    4'h5: pe14_in03 <= mem0517;
    4'h6: pe14_in03 <= mem0617;
    4'h7: pe14_in03 <= mem0717;
    4'h8: pe14_in03 <= mem0817;
    4'h9: pe14_in03 <= mem0917;
    4'ha: pe14_in03 <= mem1017;
    4'hb: pe14_in03 <= mem1117;
    4'hc: pe14_in03 <= mem1217;
    4'hd: pe14_in03 <= mem1317;
    4'he: pe14_in03 <= mem1417;
    4'hf: pe14_in03 <= mem1517;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in04 <= mem0114;
    4'h1: pe14_in04 <= mem0214;
    4'h2: pe14_in04 <= mem0314;
    4'h3: pe14_in04 <= mem0414;
    4'h4: pe14_in04 <= mem0514;
    4'h5: pe14_in04 <= mem0614;
    4'h6: pe14_in04 <= mem0714;
    4'h7: pe14_in04 <= mem0814;
    4'h8: pe14_in04 <= mem0914;
    4'h9: pe14_in04 <= mem1014;
    4'ha: pe14_in04 <= mem1114;
    4'hb: pe14_in04 <= mem1214;
    4'hc: pe14_in04 <= mem1314;
    4'hd: pe14_in04 <= mem1414;
    4'he: pe14_in04 <= mem1514;
    4'hf: pe14_in04 <= mem1614;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in05 <= mem0115;
    4'h1: pe14_in05 <= mem0215;
    4'h2: pe14_in05 <= mem0315;
    4'h3: pe14_in05 <= mem0415;
    4'h4: pe14_in05 <= mem0515;
    4'h5: pe14_in05 <= mem0615;
    4'h6: pe14_in05 <= mem0715;
    4'h7: pe14_in05 <= mem0815;
    4'h8: pe14_in05 <= mem0915;
    4'h9: pe14_in05 <= mem1015;
    4'ha: pe14_in05 <= mem1115;
    4'hb: pe14_in05 <= mem1215;
    4'hc: pe14_in05 <= mem1315;
    4'hd: pe14_in05 <= mem1415;
    4'he: pe14_in05 <= mem1515;
    4'hf: pe14_in05 <= mem1615;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in06 <= mem0116;
    4'h1: pe14_in06 <= mem0216;
    4'h2: pe14_in06 <= mem0316;
    4'h3: pe14_in06 <= mem0416;
    4'h4: pe14_in06 <= mem0516;
    4'h5: pe14_in06 <= mem0616;
    4'h6: pe14_in06 <= mem0716;
    4'h7: pe14_in06 <= mem0816;
    4'h8: pe14_in06 <= mem0916;
    4'h9: pe14_in06 <= mem1016;
    4'ha: pe14_in06 <= mem1116;
    4'hb: pe14_in06 <= mem1216;
    4'hc: pe14_in06 <= mem1316;
    4'hd: pe14_in06 <= mem1416;
    4'he: pe14_in06 <= mem1516;
    4'hf: pe14_in06 <= mem1616;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in07 <= mem0117;
    4'h1: pe14_in07 <= mem0217;
    4'h2: pe14_in07 <= mem0317;
    4'h3: pe14_in07 <= mem0417;
    4'h4: pe14_in07 <= mem0517;
    4'h5: pe14_in07 <= mem0617;
    4'h6: pe14_in07 <= mem0717;
    4'h7: pe14_in07 <= mem0817;
    4'h8: pe14_in07 <= mem0917;
    4'h9: pe14_in07 <= mem1017;
    4'ha: pe14_in07 <= mem1117;
    4'hb: pe14_in07 <= mem1217;
    4'hc: pe14_in07 <= mem1317;
    4'hd: pe14_in07 <= mem1417;
    4'he: pe14_in07 <= mem1517;
    4'hf: pe14_in07 <= mem1617;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in08 <= mem0214;
    4'h1: pe14_in08 <= mem0314;
    4'h2: pe14_in08 <= mem0414;
    4'h3: pe14_in08 <= mem0514;
    4'h4: pe14_in08 <= mem0614;
    4'h5: pe14_in08 <= mem0714;
    4'h6: pe14_in08 <= mem0814;
    4'h7: pe14_in08 <= mem0914;
    4'h8: pe14_in08 <= mem1014;
    4'h9: pe14_in08 <= mem1114;
    4'ha: pe14_in08 <= mem1214;
    4'hb: pe14_in08 <= mem1314;
    4'hc: pe14_in08 <= mem1414;
    4'hd: pe14_in08 <= mem1514;
    4'he: pe14_in08 <= mem1614;
    4'hf: pe14_in08 <= mem1714;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in09 <= mem0215;
    4'h1: pe14_in09 <= mem0315;
    4'h2: pe14_in09 <= mem0415;
    4'h3: pe14_in09 <= mem0515;
    4'h4: pe14_in09 <= mem0615;
    4'h5: pe14_in09 <= mem0715;
    4'h6: pe14_in09 <= mem0815;
    4'h7: pe14_in09 <= mem0915;
    4'h8: pe14_in09 <= mem1015;
    4'h9: pe14_in09 <= mem1115;
    4'ha: pe14_in09 <= mem1215;
    4'hb: pe14_in09 <= mem1315;
    4'hc: pe14_in09 <= mem1415;
    4'hd: pe14_in09 <= mem1515;
    4'he: pe14_in09 <= mem1615;
    4'hf: pe14_in09 <= mem1715;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in10 <= mem0216;
    4'h1: pe14_in10 <= mem0316;
    4'h2: pe14_in10 <= mem0416;
    4'h3: pe14_in10 <= mem0516;
    4'h4: pe14_in10 <= mem0616;
    4'h5: pe14_in10 <= mem0716;
    4'h6: pe14_in10 <= mem0816;
    4'h7: pe14_in10 <= mem0916;
    4'h8: pe14_in10 <= mem1016;
    4'h9: pe14_in10 <= mem1116;
    4'ha: pe14_in10 <= mem1216;
    4'hb: pe14_in10 <= mem1316;
    4'hc: pe14_in10 <= mem1416;
    4'hd: pe14_in10 <= mem1516;
    4'he: pe14_in10 <= mem1616;
    4'hf: pe14_in10 <= mem1716;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in11 <= mem0217;
    4'h1: pe14_in11 <= mem0317;
    4'h2: pe14_in11 <= mem0417;
    4'h3: pe14_in11 <= mem0517;
    4'h4: pe14_in11 <= mem0617;
    4'h5: pe14_in11 <= mem0717;
    4'h6: pe14_in11 <= mem0817;
    4'h7: pe14_in11 <= mem0917;
    4'h8: pe14_in11 <= mem1017;
    4'h9: pe14_in11 <= mem1117;
    4'ha: pe14_in11 <= mem1217;
    4'hb: pe14_in11 <= mem1317;
    4'hc: pe14_in11 <= mem1417;
    4'hd: pe14_in11 <= mem1517;
    4'he: pe14_in11 <= mem1617;
    4'hf: pe14_in11 <= mem1717;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in12 <= mem0314;
    4'h1: pe14_in12 <= mem0414;
    4'h2: pe14_in12 <= mem0514;
    4'h3: pe14_in12 <= mem0614;
    4'h4: pe14_in12 <= mem0714;
    4'h5: pe14_in12 <= mem0814;
    4'h6: pe14_in12 <= mem0914;
    4'h7: pe14_in12 <= mem1014;
    4'h8: pe14_in12 <= mem1114;
    4'h9: pe14_in12 <= mem1214;
    4'ha: pe14_in12 <= mem1314;
    4'hb: pe14_in12 <= mem1414;
    4'hc: pe14_in12 <= mem1514;
    4'hd: pe14_in12 <= mem1614;
    4'he: pe14_in12 <= mem1714;
    4'hf: pe14_in12 <= mem1814;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in13 <= mem0315;
    4'h1: pe14_in13 <= mem0415;
    4'h2: pe14_in13 <= mem0515;
    4'h3: pe14_in13 <= mem0615;
    4'h4: pe14_in13 <= mem0715;
    4'h5: pe14_in13 <= mem0815;
    4'h6: pe14_in13 <= mem0915;
    4'h7: pe14_in13 <= mem1015;
    4'h8: pe14_in13 <= mem1115;
    4'h9: pe14_in13 <= mem1215;
    4'ha: pe14_in13 <= mem1315;
    4'hb: pe14_in13 <= mem1415;
    4'hc: pe14_in13 <= mem1515;
    4'hd: pe14_in13 <= mem1615;
    4'he: pe14_in13 <= mem1715;
    4'hf: pe14_in13 <= mem1815;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in14 <= mem0316;
    4'h1: pe14_in14 <= mem0416;
    4'h2: pe14_in14 <= mem0516;
    4'h3: pe14_in14 <= mem0616;
    4'h4: pe14_in14 <= mem0716;
    4'h5: pe14_in14 <= mem0816;
    4'h6: pe14_in14 <= mem0916;
    4'h7: pe14_in14 <= mem1016;
    4'h8: pe14_in14 <= mem1116;
    4'h9: pe14_in14 <= mem1216;
    4'ha: pe14_in14 <= mem1316;
    4'hb: pe14_in14 <= mem1416;
    4'hc: pe14_in14 <= mem1516;
    4'hd: pe14_in14 <= mem1616;
    4'he: pe14_in14 <= mem1716;
    4'hf: pe14_in14 <= mem1816;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe14_in15 <= mem0317;
    4'h1: pe14_in15 <= mem0417;
    4'h2: pe14_in15 <= mem0517;
    4'h3: pe14_in15 <= mem0617;
    4'h4: pe14_in15 <= mem0717;
    4'h5: pe14_in15 <= mem0817;
    4'h6: pe14_in15 <= mem0917;
    4'h7: pe14_in15 <= mem1017;
    4'h8: pe14_in15 <= mem1117;
    4'h9: pe14_in15 <= mem1217;
    4'ha: pe14_in15 <= mem1317;
    4'hb: pe14_in15 <= mem1417;
    4'hc: pe14_in15 <= mem1517;
    4'hd: pe14_in15 <= mem1617;
    4'he: pe14_in15 <= mem1717;
    4'hf: pe14_in15 <= mem1817;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in00 <= mem0015;
    4'h1: pe15_in00 <= mem0115;
    4'h2: pe15_in00 <= mem0215;
    4'h3: pe15_in00 <= mem0315;
    4'h4: pe15_in00 <= mem0415;
    4'h5: pe15_in00 <= mem0515;
    4'h6: pe15_in00 <= mem0615;
    4'h7: pe15_in00 <= mem0715;
    4'h8: pe15_in00 <= mem0815;
    4'h9: pe15_in00 <= mem0915;
    4'ha: pe15_in00 <= mem1015;
    4'hb: pe15_in00 <= mem1115;
    4'hc: pe15_in00 <= mem1215;
    4'hd: pe15_in00 <= mem1315;
    4'he: pe15_in00 <= mem1415;
    4'hf: pe15_in00 <= mem1515;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in01 <= mem0016;
    4'h1: pe15_in01 <= mem0116;
    4'h2: pe15_in01 <= mem0216;
    4'h3: pe15_in01 <= mem0316;
    4'h4: pe15_in01 <= mem0416;
    4'h5: pe15_in01 <= mem0516;
    4'h6: pe15_in01 <= mem0616;
    4'h7: pe15_in01 <= mem0716;
    4'h8: pe15_in01 <= mem0816;
    4'h9: pe15_in01 <= mem0916;
    4'ha: pe15_in01 <= mem1016;
    4'hb: pe15_in01 <= mem1116;
    4'hc: pe15_in01 <= mem1216;
    4'hd: pe15_in01 <= mem1316;
    4'he: pe15_in01 <= mem1416;
    4'hf: pe15_in01 <= mem1516;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in02 <= mem0017;
    4'h1: pe15_in02 <= mem0117;
    4'h2: pe15_in02 <= mem0217;
    4'h3: pe15_in02 <= mem0317;
    4'h4: pe15_in02 <= mem0417;
    4'h5: pe15_in02 <= mem0517;
    4'h6: pe15_in02 <= mem0617;
    4'h7: pe15_in02 <= mem0717;
    4'h8: pe15_in02 <= mem0817;
    4'h9: pe15_in02 <= mem0917;
    4'ha: pe15_in02 <= mem1017;
    4'hb: pe15_in02 <= mem1117;
    4'hc: pe15_in02 <= mem1217;
    4'hd: pe15_in02 <= mem1317;
    4'he: pe15_in02 <= mem1417;
    4'hf: pe15_in02 <= mem1517;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in03 <= mem0018;
    4'h1: pe15_in03 <= mem0118;
    4'h2: pe15_in03 <= mem0218;
    4'h3: pe15_in03 <= mem0318;
    4'h4: pe15_in03 <= mem0418;
    4'h5: pe15_in03 <= mem0518;
    4'h6: pe15_in03 <= mem0618;
    4'h7: pe15_in03 <= mem0718;
    4'h8: pe15_in03 <= mem0818;
    4'h9: pe15_in03 <= mem0918;
    4'ha: pe15_in03 <= mem1018;
    4'hb: pe15_in03 <= mem1118;
    4'hc: pe15_in03 <= mem1218;
    4'hd: pe15_in03 <= mem1318;
    4'he: pe15_in03 <= mem1418;
    4'hf: pe15_in03 <= mem1518;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in04 <= mem0115;
    4'h1: pe15_in04 <= mem0215;
    4'h2: pe15_in04 <= mem0315;
    4'h3: pe15_in04 <= mem0415;
    4'h4: pe15_in04 <= mem0515;
    4'h5: pe15_in04 <= mem0615;
    4'h6: pe15_in04 <= mem0715;
    4'h7: pe15_in04 <= mem0815;
    4'h8: pe15_in04 <= mem0915;
    4'h9: pe15_in04 <= mem1015;
    4'ha: pe15_in04 <= mem1115;
    4'hb: pe15_in04 <= mem1215;
    4'hc: pe15_in04 <= mem1315;
    4'hd: pe15_in04 <= mem1415;
    4'he: pe15_in04 <= mem1515;
    4'hf: pe15_in04 <= mem1615;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in05 <= mem0116;
    4'h1: pe15_in05 <= mem0216;
    4'h2: pe15_in05 <= mem0316;
    4'h3: pe15_in05 <= mem0416;
    4'h4: pe15_in05 <= mem0516;
    4'h5: pe15_in05 <= mem0616;
    4'h6: pe15_in05 <= mem0716;
    4'h7: pe15_in05 <= mem0816;
    4'h8: pe15_in05 <= mem0916;
    4'h9: pe15_in05 <= mem1016;
    4'ha: pe15_in05 <= mem1116;
    4'hb: pe15_in05 <= mem1216;
    4'hc: pe15_in05 <= mem1316;
    4'hd: pe15_in05 <= mem1416;
    4'he: pe15_in05 <= mem1516;
    4'hf: pe15_in05 <= mem1616;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in06 <= mem0117;
    4'h1: pe15_in06 <= mem0217;
    4'h2: pe15_in06 <= mem0317;
    4'h3: pe15_in06 <= mem0417;
    4'h4: pe15_in06 <= mem0517;
    4'h5: pe15_in06 <= mem0617;
    4'h6: pe15_in06 <= mem0717;
    4'h7: pe15_in06 <= mem0817;
    4'h8: pe15_in06 <= mem0917;
    4'h9: pe15_in06 <= mem1017;
    4'ha: pe15_in06 <= mem1117;
    4'hb: pe15_in06 <= mem1217;
    4'hc: pe15_in06 <= mem1317;
    4'hd: pe15_in06 <= mem1417;
    4'he: pe15_in06 <= mem1517;
    4'hf: pe15_in06 <= mem1617;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in07 <= mem0118;
    4'h1: pe15_in07 <= mem0218;
    4'h2: pe15_in07 <= mem0318;
    4'h3: pe15_in07 <= mem0418;
    4'h4: pe15_in07 <= mem0518;
    4'h5: pe15_in07 <= mem0618;
    4'h6: pe15_in07 <= mem0718;
    4'h7: pe15_in07 <= mem0818;
    4'h8: pe15_in07 <= mem0918;
    4'h9: pe15_in07 <= mem1018;
    4'ha: pe15_in07 <= mem1118;
    4'hb: pe15_in07 <= mem1218;
    4'hc: pe15_in07 <= mem1318;
    4'hd: pe15_in07 <= mem1418;
    4'he: pe15_in07 <= mem1518;
    4'hf: pe15_in07 <= mem1618;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in08 <= mem0215;
    4'h1: pe15_in08 <= mem0315;
    4'h2: pe15_in08 <= mem0415;
    4'h3: pe15_in08 <= mem0515;
    4'h4: pe15_in08 <= mem0615;
    4'h5: pe15_in08 <= mem0715;
    4'h6: pe15_in08 <= mem0815;
    4'h7: pe15_in08 <= mem0915;
    4'h8: pe15_in08 <= mem1015;
    4'h9: pe15_in08 <= mem1115;
    4'ha: pe15_in08 <= mem1215;
    4'hb: pe15_in08 <= mem1315;
    4'hc: pe15_in08 <= mem1415;
    4'hd: pe15_in08 <= mem1515;
    4'he: pe15_in08 <= mem1615;
    4'hf: pe15_in08 <= mem1715;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in09 <= mem0216;
    4'h1: pe15_in09 <= mem0316;
    4'h2: pe15_in09 <= mem0416;
    4'h3: pe15_in09 <= mem0516;
    4'h4: pe15_in09 <= mem0616;
    4'h5: pe15_in09 <= mem0716;
    4'h6: pe15_in09 <= mem0816;
    4'h7: pe15_in09 <= mem0916;
    4'h8: pe15_in09 <= mem1016;
    4'h9: pe15_in09 <= mem1116;
    4'ha: pe15_in09 <= mem1216;
    4'hb: pe15_in09 <= mem1316;
    4'hc: pe15_in09 <= mem1416;
    4'hd: pe15_in09 <= mem1516;
    4'he: pe15_in09 <= mem1616;
    4'hf: pe15_in09 <= mem1716;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in10 <= mem0217;
    4'h1: pe15_in10 <= mem0317;
    4'h2: pe15_in10 <= mem0417;
    4'h3: pe15_in10 <= mem0517;
    4'h4: pe15_in10 <= mem0617;
    4'h5: pe15_in10 <= mem0717;
    4'h6: pe15_in10 <= mem0817;
    4'h7: pe15_in10 <= mem0917;
    4'h8: pe15_in10 <= mem1017;
    4'h9: pe15_in10 <= mem1117;
    4'ha: pe15_in10 <= mem1217;
    4'hb: pe15_in10 <= mem1317;
    4'hc: pe15_in10 <= mem1417;
    4'hd: pe15_in10 <= mem1517;
    4'he: pe15_in10 <= mem1617;
    4'hf: pe15_in10 <= mem1717;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in11 <= mem0218;
    4'h1: pe15_in11 <= mem0318;
    4'h2: pe15_in11 <= mem0418;
    4'h3: pe15_in11 <= mem0518;
    4'h4: pe15_in11 <= mem0618;
    4'h5: pe15_in11 <= mem0718;
    4'h6: pe15_in11 <= mem0818;
    4'h7: pe15_in11 <= mem0918;
    4'h8: pe15_in11 <= mem1018;
    4'h9: pe15_in11 <= mem1118;
    4'ha: pe15_in11 <= mem1218;
    4'hb: pe15_in11 <= mem1318;
    4'hc: pe15_in11 <= mem1418;
    4'hd: pe15_in11 <= mem1518;
    4'he: pe15_in11 <= mem1618;
    4'hf: pe15_in11 <= mem1718;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in12 <= mem0315;
    4'h1: pe15_in12 <= mem0415;
    4'h2: pe15_in12 <= mem0515;
    4'h3: pe15_in12 <= mem0615;
    4'h4: pe15_in12 <= mem0715;
    4'h5: pe15_in12 <= mem0815;
    4'h6: pe15_in12 <= mem0915;
    4'h7: pe15_in12 <= mem1015;
    4'h8: pe15_in12 <= mem1115;
    4'h9: pe15_in12 <= mem1215;
    4'ha: pe15_in12 <= mem1315;
    4'hb: pe15_in12 <= mem1415;
    4'hc: pe15_in12 <= mem1515;
    4'hd: pe15_in12 <= mem1615;
    4'he: pe15_in12 <= mem1715;
    4'hf: pe15_in12 <= mem1815;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in13 <= mem0316;
    4'h1: pe15_in13 <= mem0416;
    4'h2: pe15_in13 <= mem0516;
    4'h3: pe15_in13 <= mem0616;
    4'h4: pe15_in13 <= mem0716;
    4'h5: pe15_in13 <= mem0816;
    4'h6: pe15_in13 <= mem0916;
    4'h7: pe15_in13 <= mem1016;
    4'h8: pe15_in13 <= mem1116;
    4'h9: pe15_in13 <= mem1216;
    4'ha: pe15_in13 <= mem1316;
    4'hb: pe15_in13 <= mem1416;
    4'hc: pe15_in13 <= mem1516;
    4'hd: pe15_in13 <= mem1616;
    4'he: pe15_in13 <= mem1716;
    4'hf: pe15_in13 <= mem1816;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in14 <= mem0317;
    4'h1: pe15_in14 <= mem0417;
    4'h2: pe15_in14 <= mem0517;
    4'h3: pe15_in14 <= mem0617;
    4'h4: pe15_in14 <= mem0717;
    4'h5: pe15_in14 <= mem0817;
    4'h6: pe15_in14 <= mem0917;
    4'h7: pe15_in14 <= mem1017;
    4'h8: pe15_in14 <= mem1117;
    4'h9: pe15_in14 <= mem1217;
    4'ha: pe15_in14 <= mem1317;
    4'hb: pe15_in14 <= mem1417;
    4'hc: pe15_in14 <= mem1517;
    4'hd: pe15_in14 <= mem1617;
    4'he: pe15_in14 <= mem1717;
    4'hf: pe15_in14 <= mem1817;
    endcase
end

always @ (clk)
    begin
    case (ctr_word)
    4'h0: pe15_in15 <= mem0318;
    4'h1: pe15_in15 <= mem0418;
    4'h2: pe15_in15 <= mem0518;
    4'h3: pe15_in15 <= mem0618;
    4'h4: pe15_in15 <= mem0718;
    4'h5: pe15_in15 <= mem0818;
    4'h6: pe15_in15 <= mem0918;
    4'h7: pe15_in15 <= mem1018;
    4'h8: pe15_in15 <= mem1118;
    4'h9: pe15_in15 <= mem1218;
    4'ha: pe15_in15 <= mem1318;
    4'hb: pe15_in15 <= mem1418;
    4'hc: pe15_in15 <= mem1518;
    4'hd: pe15_in15 <= mem1618;
    4'he: pe15_in15 <= mem1718;
    4'hf: pe15_in15 <= mem1818;
    endcase
end
/************************OUTPUT Logic END************************/
endmodule