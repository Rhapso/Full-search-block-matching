/**************************************************************** 
  ** Title : top module
  ** Project :  full-search block matching algorithm on VLSI
***************************************************************** 
  ** File :  top.v
  ** Author : fzp
  ** Organization: sjtu
  ** Created :  
  ** Last update : 
  ** Platform : 
  ** Simulators : 
  ** Synthesizers: 
  ** Targets : 
  ** Dependency :  
***************************************************************** 
  ** Description:  
***************************************************************** 
  ** Copyright (c) notice  
*****************************************************************/ 
module top
#(
    parameter WORD_WIDETH =                 8
)
(
    input clk,
    input en_init,
    input input_raw,
    input rst_n,
    output reg serial20
);

endmodule